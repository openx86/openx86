/*
project: w80386dx
author: Chang Wei<changwei1006@gmail.com>
repo: https://github.com/openx86/w80386dx
module: decode unit
create at: 2022-01-04 03:27:51
description: decode unit module
*/

`include "D:/GitHub/openx86/w80386dx/rtl/definition.h"

module decode (
    input  logic [ 7:0] i_instruction [0:15],
    input  logic        i_default_operand_size,
    output logic        o_opcode_x86_AAA_ASCII_adjust_after_add,
    output logic        o_opcode_x86_AAD_ASCII_AX_before_div,
    output logic        o_opcode_x86_AAM_ASCII_AX_after_mul,
    output logic        o_opcode_x86_AAS_ASCII_adjust_after_sub,
    output logic        o_opcode_x86_ADC_reg_to_reg_mem,
    output logic        o_opcode_x86_ADC_reg_mem_to_reg,
    output logic        o_opcode_x86_ADC_imm_to_reg_mem,
    output logic        o_opcode_x86_ADC_imm_to_acc,
    output logic        o_opcode_x86_ADD_reg_to_reg_mem,
    output logic        o_opcode_x86_ADD_reg_mem_to_reg,
    output logic        o_opcode_x86_ADD_imm_to_reg_mem,
    output logic        o_opcode_x86_ADD_imm_to_acc,
    output logic        o_opcode_x86_AND_reg_to_reg_mem,
    output logic        o_opcode_x86_AND_reg_mem_to_reg,
    output logic        o_opcode_x86_AND_imm_to_reg_mem,
    output logic        o_opcode_x86_AND_imm_to_acc,
    output logic        o_opcode_x86_ARPL_adjust_RPL_field_of_selector,
    output logic        o_opcode_x86_BOUND_check_array_against_bounds,
    output logic        o_opcode_x86_BSF_bit_scan_forward,
    output logic        o_opcode_x86_BSR_bit_scan_reverse,
    output logic        o_opcode_x86_BSWAP_byte_swap,
    output logic        o_opcode_x86_BT_reg_mem_with_imm,
    output logic        o_opcode_x86_BT_reg_mem_with_reg,
    output logic        o_opcode_x86_BTC_reg_mem_with_imm,
    output logic        o_opcode_x86_BTC_reg_mem_with_reg,
    output logic        o_opcode_x86_BTR_reg_mem_with_imm,
    output logic        o_opcode_x86_BTR_reg_mem_with_reg,
    output logic        o_opcode_x86_BTS_reg_mem_with_imm,
    output logic        o_opcode_x86_BTS_reg_mem_with_reg,
    output logic        o_opcode_x86_CALL_in_same_segment_direct,
    output logic        o_opcode_x86_CALL_in_same_segment_indirec,
    output logic        o_opcode_x86_CALL_in_other_segment_direct,
    output logic        o_opcode_x86_CALL_in_other_segment_indirect,
    output logic        o_opcode_x86_CBW_convert_byte_to_word,
    output logic        o_opcode_x86_CDQ_convert_double_word_to_quad_word,
    output logic        o_opcode_x86_CLC_clear_carry_flag,
    output logic        o_opcode_x86_CLD_clear_direction_flag,
    output logic        o_opcode_x86_CLI_clear_interrupt_enable_flag,
    output logic        o_opcode_x86_CLTS_clear_task_switched_flag,
    output logic        o_opcode_x86_CMC_complement_carry_flag,
    output logic        o_opcode_x86_CMP_mem_with_reg,
    output logic        o_opcode_x86_CMP_reg_with_mem,
    output logic        o_opcode_x86_CMP_imm_with_reg_mem,
    output logic        o_opcode_x86_CMP_imm_with_acc,
    output logic        o_opcode_x86_CMPS_compare_string_operands,
    output logic        o_opcode_x86_CMPXCHG_compare_and_exchange,
    output logic        o_opcode_x86_CPUID_CPU_identification,
    output logic        o_opcode_x86_CWD_convert_word_to_double,
    output logic        o_opcode_x86_CWDE_convert_word_to_double,
    output logic        o_opcode_x86_DAA_decimal_adjust_AL_after_add,
    output logic        o_opcode_x86_DAS_decimal_adjust_AL_after_sub,
    output logic        o_opcode_x86_DEC_reg_mem,
    output logic        o_opcode_x86_DEC_reg,
    output logic        o_opcode_x86_DIV_acc_by_reg_mem,
    output logic        o_opcode_x86_HLT_halt,
    output logic        o_opcode_x86_IDIV_acc_by_reg_mem,
    output logic        o_opcode_x86_IMUL_acc_with_reg_mem,
    output logic        o_opcode_x86_IMUL_reg_with_reg_mem,
    output logic        o_opcode_x86_IMUL_reg_mem_with_imm_to_reg,
    output logic        o_opcode_x86_IN_port_fixed,
    output logic        o_opcode_x86_IN_port_variable,
    output logic        o_opcode_x86_INC_reg_mem,
    output logic        o_opcode_x86_INC_reg,
    output logic        o_opcode_x86_INS_input_from_DX_port,
    output logic        o_opcode_x86_INT_interrupt_type_n,
    output logic        o_opcode_x86_INT_interrupt_type_3,
    output logic        o_opcode_x86_INT_interrupt_type_4,
    output logic        o_opcode_x86_INVD_invalidate_cache,
    output logic        o_opcode_x86_INVLPG_invalidate_TLB_entry,
    output logic        o_opcode_x86_INVPCID_invalidate_process_ctx_id,
    output logic        o_opcode_x86_IRET_interrupt_return,
    output logic        o_opcode_x86_Jcc_jump_if_cond_is_met_8_bit_disp,
    output logic        o_opcode_x86_Jcc_jump_if_cond_is_met_full_disp,
    output logic        o_opcode_x86_JCXZ_jump_on_CX_zero,
    output logic        o_opcode_x86_JMP_to_same_segment_short,
    output logic        o_opcode_x86_JMP_to_same_segment_direct,
    output logic        o_opcode_x86_JMP_to_same_segment_indirect,
    output logic        o_opcode_x86_JMP_to_other_segment_direct,
    output logic        o_opcode_x86_JMP_to_other_segment_indirect,
    output logic        o_opcode_x86_LAHF_load_FLAG_into_AH,
    output logic        o_opcode_x86_LAR_load_access_rights_byte,
    output logic        o_opcode_x86_LDS_load_pointer_to_DS,
    output logic        o_opcode_x86_LEA_load_effective_adddress_to_reg,
    output logic        o_opcode_x86_LEAVE_high_level_procedure_exit,
    output logic        o_opcode_x86_LES_load_pointer_to_ES,
    output logic        o_opcode_x86_LFS_load_pointer_to_FS,
    output logic        o_opcode_x86_LGDT_load_global_desciptor_table_reg,
    output logic        o_opcode_x86_LGS_load_pointer_to_GS,
    output logic        o_opcode_x86_LIDT_load_interrupt_desciptor_table_reg,
    output logic        o_opcode_x86_LLDT_load_local_desciptor_table_reg,
    output logic        o_opcode_x86_LMSW_load_status_word,
    output logic        o_opcode_x86_LODS_load_string_operand,
    output logic        o_opcode_x86_LOOP_count,
    output logic        o_opcode_x86_LOOPZ_count_while_zero,
    output logic        o_opcode_x86_LOOPNZ_count_while_not_zero,
    output logic        o_opcode_x86_LSL_load_segment_limit,
    output logic        o_opcode_x86_LSS_load_pointer_to_SS,
    output logic        o_opcode_x86_LTR_load_task_register,
    output logic        o_opcode_x86_MOV_reg_to_reg_mem,
    output logic        o_opcode_x86_MOV_reg_mem_to_reg,
    output logic        o_opcode_x86_MOV_imm_to_reg_mem,
    output logic        o_opcode_x86_MOV_imm_to_reg,
    output logic        o_opcode_x86_MOV_mem_to_acc,
    output logic        o_opcode_x86_MOV_acc_to_mem,
    output logic        o_opcode_x86_MOV_CR_from_reg,
    output logic        o_opcode_x86_MOV_reg_from_CR,
    output logic        o_opcode_x86_MOV_DR_from_reg,
    output logic        o_opcode_x86_MOV_reg_from_DR,
    output logic        o_opcode_x86_MOV_TR_from_reg,
    output logic        o_opcode_x86_MOV_reg_from_TR,
    output logic        o_opcode_x86_MOV_reg_mem_to_sreg,
    output logic        o_opcode_x86_MOV_sreg_to_reg_mem,
    output logic        o_opcode_x86_MOVBE_move_data_after_swapping_bytes_reg_mem_to_reg,
    output logic        o_opcode_x86_MOVBE_move_data_after_swapping_bytes_reg_to_reg_mem,
    output logic        o_opcode_x86_MOVS_move_data_from_string_to_string,
    output logic        o_opcode_x86_MOVSX_move_with_sign_extend_mem_reg_to_reg,
    output logic        o_opcode_x86_MOVZX_move_with_zero_extend_mem_reg_to_reg,
    output logic        o_opcode_x86_MUL_acc_with_reg_mem,
    output logic        o_opcode_x86_NEG_two_s_complement_negation,
    output logic        o_opcode_x86_NOP_no_operation,
    output logic        o_opcode_x86_NOP_no_operation_multi_byte,
    output logic        o_opcode_x86_NOT_one_s_complement_negation,
    output logic        o_opcode_x86_OR_reg_to_reg_mem,
    output logic        o_opcode_x86_OR_reg_mem_to_reg,
    output logic        o_opcode_x86_OR_imm_to_reg_mem,
    output logic        o_opcode_x86_OR_imm_to_acc,
    output logic        o_opcode_x86_OUT_port_fixed,
    output logic        o_opcode_x86_OUT_port_variable,
    output logic        o_opcode_x86_OUTS_output_string,
    output logic        o_opcode_x86_POP_reg_mem,
    output logic        o_opcode_x86_POP_reg,
    output logic        o_opcode_x86_POP_sreg_2,
    output logic        o_opcode_x86_POP_sreg_3,
    output logic        o_opcode_x86_POPA_pop_all_general_registers,
    output logic        o_opcode_x86_POPF_pop_stack_into_FLAGS_or_EFLAGS,
    output logic        o_opcode_x86_PUSH_reg_mem,
    output logic        o_opcode_x86_PUSH_reg,
    output logic        o_opcode_x86_PUSH_sreg_2,
    output logic        o_opcode_x86_PUSH_sreg_3,
    output logic        o_opcode_x86_PUSH_imm,
    output logic        o_opcode_x86_PUSH_all_general_registers,
    output logic        o_opcode_x86_PUSHF_push_flags_onto_stack,
    output logic        o_opcode_x86_RCL_reg_mem_by_1,
    output logic        o_opcode_x86_RCL_reg_mem_by_CL,
    output logic        o_opcode_x86_RCL_reg_mem_by_imm,
    output logic        o_opcode_x86_RCR_reg_mem_by_1,
    output logic        o_opcode_x86_RCR_reg_mem_by_CL,
    output logic        o_opcode_x86_RCR_reg_mem_by_imm,
    output logic        o_opcode_x86_RDMSR_read_from_model_specific_reg,
    output logic        o_opcode_x86_RDPCM_read_performance_monitoring_counters,
    output logic        o_opcode_x86_RDTSC_read_time_stamp_counter,
    output logic        o_opcode_x86_RDTSC_read_time_stamp_counter_and_processor_id,
    output logic        o_opcode_x86_REP_INS_input_string,
    output logic        o_opcode_x86_REP_LODS_load_string,
    output logic        o_opcode_x86_REP_MOVS_move_string,
    output logic        o_opcode_x86_REP_OUTS_output_string,
    output logic        o_opcode_x86_REP_STOS_store_string,
    output logic        o_opcode_x86_REPE_CMPS_compare_string,
    output logic        o_opcode_x86_REPE_SCAS_scan_string,
    output logic        o_opcode_x86_REPNE_CMPS_compare_string,
    output logic        o_opcode_x86_REPNE_SCAS_scan_string,
    output logic        o_opcode_x86_RET_return_from_procedure_to_same_segment_no_argument,
    output logic        o_opcode_x86_RET_return_from_procedure_to_same_segment_adding_imm_to_SP,
    output logic        o_opcode_x86_RET_return_from_procedure_to_other_segment_no_argument,
    output logic        o_opcode_x86_RET_return_from_procedure_to_other_segment_adding_imm_to_SP,
    output logic        o_opcode_x86_ROL_reg_mem_by_1,
    output logic        o_opcode_x86_ROL_reg_mem_by_CL,
    output logic        o_opcode_x86_ROL_reg_mem_by_imm,
    output logic        o_opcode_x86_ROR_reg_mem_by_1,
    output logic        o_opcode_x86_ROR_reg_mem_by_CL,
    output logic        o_opcode_x86_ROR_reg_mem_by_imm,
    output logic        o_opcode_x86_RSM_resume_from_system_management_mode,
    output logic        o_opcode_x86_SAHF_store_AH_into_flags,
    output logic        o_opcode_x86_SAR_reg_mem_by_1,
    output logic        o_opcode_x86_SAR_reg_mem_by_CL,
    output logic        o_opcode_x86_SAR_reg_mem_by_imm,
    output logic        o_opcode_x86_SBB_reg_to_reg_mem,
    output logic        o_opcode_x86_SBB_reg_mem_to_reg,
    output logic        o_opcode_x86_SBB_imm_to_reg_mem,
    output logic        o_opcode_x86_SBB_imm_to_acc,
    output logic        o_opcode_x86_SCAS_scan_string,
    output logic        o_opcode_x86_SETcc_byte_set_on_condition,
    output logic        o_opcode_x86_SGDT_store_global_descriptor_table_register,
    output logic        o_opcode_x86_SHL_reg_mem_by_1,
    output logic        o_opcode_x86_SHL_reg_mem_by_CL,
    output logic        o_opcode_x86_SHL_reg_mem_by_imm,
    output logic        o_opcode_x86_SHLD_reg_mem_by_imm,
    output logic        o_opcode_x86_SHLD_reg_mem_by_CL,
    output logic        o_opcode_x86_SHR_reg_mem_by_1,
    output logic        o_opcode_x86_SHR_reg_mem_by_CL,
    output logic        o_opcode_x86_SHR_reg_mem_by_imm,
    output logic        o_opcode_x86_SHRD_reg_mem_by_imm,
    output logic        o_opcode_x86_SHRD_reg_mem_by_CL,
    output logic        o_opcode_x86_SIDT_store_interrupt_desciptor_table_register,
    output logic        o_opcode_x86_SLDT_store_local_desciptor_table_register,
    output logic        o_opcode_x86_SMSW_store_machine_status_word,
    output logic        o_opcode_x86_STC_set_carry_flag,
    output logic        o_opcode_x86_STD_set_direction_flag,
    output logic        o_opcode_x86_STI_set_interrupt_enable_flag,
    output logic        o_opcode_x86_STOS_store_string_data,
    output logic        o_opcode_x86_STR_store_task_register,
    output logic        o_opcode_x86_SUB_reg_to_reg_mem,
    output logic        o_opcode_x86_SUB_reg_mem_to_reg,
    output logic        o_opcode_x86_SUB_imm_to_reg_mem,
    output logic        o_opcode_x86_SUB_imm_to_acc,
    output logic        o_opcode_x86_TEST_reg_mem_and_reg,
    output logic        o_opcode_x86_TEST_imm_and_reg_mem,
    output logic        o_opcode_x86_TEST_imm_and_acc,
    output logic        o_opcode_x86_UD0_undefined_instruction,
    output logic        o_opcode_x86_UD1_undefined_instruction,
    output logic        o_opcode_x86_UD2_undefined_instruction,
    output logic        o_opcode_x86_VERR_verify_a_segment_for_reading,
    output logic        o_opcode_x86_VERW_verify_a_segment_for_writing,
    output logic        o_opcode_x86_WAIT_wait,
    output logic        o_opcode_x86_WBINVD_writeback_and_invalidate_data_cache,
    output logic        o_opcode_x86_WRMSR_write_to_model_specific_register,
    output logic        o_opcode_x86_XADD_exchange_and_add,
    output logic        o_opcode_x86_XCHG_reg_mem_with_reg,
    output logic        o_opcode_x86_XCHG_reg_with_acc_short,
    output logic        o_opcode_x86_XLAT_table_look_up_translation,
    output logic        o_opcode_x86_XOR_reg_to_reg_mem,
    output logic        o_opcode_x86_XOR_reg_mem_to_reg,
    output logic        o_opcode_x86_XOR_imm_to_reg_mem,
    output logic        o_opcode_x86_XOR_imm_to_acc,
    output logic        o_error
);

decode_opcode_x86 (
    .o_opcode_x86_AAA_ASCII_adjust_after_add ( o_opcode_x86_AAA_ASCII_adjust_after_add ),
    .o_opcode_x86_AAD_ASCII_AX_before_div ( o_opcode_x86_AAD_ASCII_AX_before_div ),
    .o_opcode_x86_AAM_ASCII_AX_after_mul ( o_opcode_x86_AAM_ASCII_AX_after_mul ),
    .o_opcode_x86_AAS_ASCII_adjust_after_sub ( o_opcode_x86_AAS_ASCII_adjust_after_sub ),
    .o_opcode_x86_ADC_reg_to_reg_mem ( o_opcode_x86_ADC_reg_to_reg_mem ),
    .o_opcode_x86_ADC_reg_mem_to_reg ( o_opcode_x86_ADC_reg_mem_to_reg ),
    .o_opcode_x86_ADC_imm_to_reg_mem ( o_opcode_x86_ADC_imm_to_reg_mem ),
    .o_opcode_x86_ADC_imm_to_acc ( o_opcode_x86_ADC_imm_to_acc ),
    .o_opcode_x86_ADD_reg_to_reg_mem ( o_opcode_x86_ADD_reg_to_reg_mem ),
    .o_opcode_x86_ADD_reg_mem_to_reg ( o_opcode_x86_ADD_reg_mem_to_reg ),
    .o_opcode_x86_ADD_imm_to_reg_mem ( o_opcode_x86_ADD_imm_to_reg_mem ),
    .o_opcode_x86_ADD_imm_to_acc ( o_opcode_x86_ADD_imm_to_acc ),
    .o_opcode_x86_AND_reg_to_reg_mem ( o_opcode_x86_AND_reg_to_reg_mem ),
    .o_opcode_x86_AND_reg_mem_to_reg ( o_opcode_x86_AND_reg_mem_to_reg ),
    .o_opcode_x86_AND_imm_to_reg_mem ( o_opcode_x86_AND_imm_to_reg_mem ),
    .o_opcode_x86_AND_imm_to_acc ( o_opcode_x86_AND_imm_to_acc ),
    .o_opcode_x86_ARPL_adjust_RPL_field_of_selector ( o_opcode_x86_ARPL_adjust_RPL_field_of_selector ),
    .o_opcode_x86_BOUND_check_array_against_bounds ( o_opcode_x86_BOUND_check_array_against_bounds ),
    .o_opcode_x86_BSF_bit_scan_forward ( o_opcode_x86_BSF_bit_scan_forward ),
    .o_opcode_x86_BSR_bit_scan_reverse ( o_opcode_x86_BSR_bit_scan_reverse ),
    .o_opcode_x86_BSWAP_byte_swap ( o_opcode_x86_BSWAP_byte_swap ),
    .o_opcode_x86_BT_reg_mem_with_imm ( o_opcode_x86_BT_reg_mem_with_imm ),
    .o_opcode_x86_BT_reg_mem_with_reg ( o_opcode_x86_BT_reg_mem_with_reg ),
    .o_opcode_x86_BTC_reg_mem_with_imm ( o_opcode_x86_BTC_reg_mem_with_imm ),
    .o_opcode_x86_BTC_reg_mem_with_reg ( o_opcode_x86_BTC_reg_mem_with_reg ),
    .o_opcode_x86_BTR_reg_mem_with_imm ( o_opcode_x86_BTR_reg_mem_with_imm ),
    .o_opcode_x86_BTR_reg_mem_with_reg ( o_opcode_x86_BTR_reg_mem_with_reg ),
    .o_opcode_x86_BTS_reg_mem_with_imm ( o_opcode_x86_BTS_reg_mem_with_imm ),
    .o_opcode_x86_BTS_reg_mem_with_reg ( o_opcode_x86_BTS_reg_mem_with_reg ),
    .o_opcode_x86_CALL_in_same_segment_direct ( o_opcode_x86_CALL_in_same_segment_direct ),
    .o_opcode_x86_CALL_in_same_segment_indirec ( o_opcode_x86_CALL_in_same_segment_indirec ),
    .o_opcode_x86_CALL_in_other_segment_direct ( o_opcode_x86_CALL_in_other_segment_direct ),
    .o_opcode_x86_CALL_in_other_segment_indirect ( o_opcode_x86_CALL_in_other_segment_indirect ),
    .o_opcode_x86_CBW_convert_byte_to_word ( o_opcode_x86_CBW_convert_byte_to_word ),
    .o_opcode_x86_CDQ_convert_double_word_to_quad_word ( o_opcode_x86_CDQ_convert_double_word_to_quad_word ),
    .o_opcode_x86_CLC_clear_carry_flag ( o_opcode_x86_CLC_clear_carry_flag ),
    .o_opcode_x86_CLD_clear_direction_flag ( o_opcode_x86_CLD_clear_direction_flag ),
    .o_opcode_x86_CLI_clear_interrupt_enable_flag ( o_opcode_x86_CLI_clear_interrupt_enable_flag ),
    .o_opcode_x86_CLTS_clear_task_switched_flag ( o_opcode_x86_CLTS_clear_task_switched_flag ),
    .o_opcode_x86_CMC_complement_carry_flag ( o_opcode_x86_CMC_complement_carry_flag ),
    .o_opcode_x86_CMP_mem_with_reg ( o_opcode_x86_CMP_mem_with_reg ),
    .o_opcode_x86_CMP_reg_with_mem ( o_opcode_x86_CMP_reg_with_mem ),
    .o_opcode_x86_CMP_imm_with_reg_mem ( o_opcode_x86_CMP_imm_with_reg_mem ),
    .o_opcode_x86_CMP_imm_with_acc ( o_opcode_x86_CMP_imm_with_acc ),
    .o_opcode_x86_CMPS_compare_string_operands ( o_opcode_x86_CMPS_compare_string_operands ),
    .o_opcode_x86_CMPXCHG_compare_and_exchange ( o_opcode_x86_CMPXCHG_compare_and_exchange ),
    .o_opcode_x86_CPUID_CPU_identification ( o_opcode_x86_CPUID_CPU_identification ),
    .o_opcode_x86_CWD_convert_word_to_double ( o_opcode_x86_CWD_convert_word_to_double ),
    .o_opcode_x86_CWDE_convert_word_to_double ( o_opcode_x86_CWDE_convert_word_to_double ),
    .o_opcode_x86_DAA_decimal_adjust_AL_after_add ( o_opcode_x86_DAA_decimal_adjust_AL_after_add ),
    .o_opcode_x86_DAS_decimal_adjust_AL_after_sub ( o_opcode_x86_DAS_decimal_adjust_AL_after_sub ),
    .o_opcode_x86_DEC_reg_mem ( o_opcode_x86_DEC_reg_mem ),
    .o_opcode_x86_DEC_reg ( o_opcode_x86_DEC_reg ),
    .o_opcode_x86_DIV_acc_by_reg_mem ( o_opcode_x86_DIV_acc_by_reg_mem ),
    .o_opcode_x86_HLT_halt ( o_opcode_x86_HLT_halt ),
    .o_opcode_x86_IDIV_acc_by_reg_mem ( o_opcode_x86_IDIV_acc_by_reg_mem ),
    .o_opcode_x86_IMUL_acc_with_reg_mem ( o_opcode_x86_IMUL_acc_with_reg_mem ),
    .o_opcode_x86_IMUL_reg_with_reg_mem ( o_opcode_x86_IMUL_reg_with_reg_mem ),
    .o_opcode_x86_IMUL_reg_mem_with_imm_to_reg ( o_opcode_x86_IMUL_reg_mem_with_imm_to_reg ),
    .o_opcode_x86_IN_port_fixed ( o_opcode_x86_IN_port_fixed ),
    .o_opcode_x86_IN_port_variable ( o_opcode_x86_IN_port_variable ),
    .o_opcode_x86_INC_reg_mem ( o_opcode_x86_INC_reg_mem ),
    .o_opcode_x86_INC_reg ( o_opcode_x86_INC_reg ),
    .o_opcode_x86_INS_input_from_DX_port ( o_opcode_x86_INS_input_from_DX_port ),
    .o_opcode_x86_INT_interrupt_type_n ( o_opcode_x86_INT_interrupt_type_n ),
    .o_opcode_x86_INT_interrupt_type_3 ( o_opcode_x86_INT_interrupt_type_3 ),
    .o_opcode_x86_INT_interrupt_type_4 ( o_opcode_x86_INT_interrupt_type_4 ),
    .o_opcode_x86_INVD_invalidate_cache ( o_opcode_x86_INVD_invalidate_cache ),
    .o_opcode_x86_INVLPG_invalidate_TLB_entry ( o_opcode_x86_INVLPG_invalidate_TLB_entry ),
    .o_opcode_x86_INVPCID_invalidate_process_ctx_id ( o_opcode_x86_INVPCID_invalidate_process_ctx_id ),
    .o_opcode_x86_IRET_interrupt_return ( o_opcode_x86_IRET_interrupt_return ),
    .o_opcode_x86_Jcc_jump_if_cond_is_met_8_bit_disp ( o_opcode_x86_Jcc_jump_if_cond_is_met_8_bit_disp ),
    .o_opcode_x86_Jcc_jump_if_cond_is_met_full_disp ( o_opcode_x86_Jcc_jump_if_cond_is_met_full_disp ),
    .o_opcode_x86_JCXZ_jump_on_CX_zero ( o_opcode_x86_JCXZ_jump_on_CX_zero ),
    .o_opcode_x86_JMP_to_same_segment_short ( o_opcode_x86_JMP_to_same_segment_short ),
    .o_opcode_x86_JMP_to_same_segment_direct ( o_opcode_x86_JMP_to_same_segment_direct ),
    .o_opcode_x86_JMP_to_same_segment_indirect ( o_opcode_x86_JMP_to_same_segment_indirect ),
    .o_opcode_x86_JMP_to_other_segment_direct ( o_opcode_x86_JMP_to_other_segment_direct ),
    .o_opcode_x86_JMP_to_other_segment_indirect ( o_opcode_x86_JMP_to_other_segment_indirect ),
    .o_opcode_x86_LAHF_load_FLAG_into_AH ( o_opcode_x86_LAHF_load_FLAG_into_AH ),
    .o_opcode_x86_LAR_load_access_rights_byte ( o_opcode_x86_LAR_load_access_rights_byte ),
    .o_opcode_x86_LDS_load_pointer_to_DS ( o_opcode_x86_LDS_load_pointer_to_DS ),
    .o_opcode_x86_LEA_load_effective_adddress_to_reg ( o_opcode_x86_LEA_load_effective_adddress_to_reg ),
    .o_opcode_x86_LEAVE_high_level_procedure_exit ( o_opcode_x86_LEAVE_high_level_procedure_exit ),
    .o_opcode_x86_LES_load_pointer_to_ES ( o_opcode_x86_LES_load_pointer_to_ES ),
    .o_opcode_x86_LFS_load_pointer_to_FS ( o_opcode_x86_LFS_load_pointer_to_FS ),
    .o_opcode_x86_LGDT_load_global_desciptor_table_reg ( o_opcode_x86_LGDT_load_global_desciptor_table_reg ),
    .o_opcode_x86_LGS_load_pointer_to_GS ( o_opcode_x86_LGS_load_pointer_to_GS ),
    .o_opcode_x86_LIDT_load_interrupt_desciptor_table_reg ( o_opcode_x86_LIDT_load_interrupt_desciptor_table_reg ),
    .o_opcode_x86_LLDT_load_local_desciptor_table_reg ( o_opcode_x86_LLDT_load_local_desciptor_table_reg ),
    .o_opcode_x86_LMSW_load_status_word ( o_opcode_x86_LMSW_load_status_word ),
    .o_opcode_x86_LODS_load_string_operand ( o_opcode_x86_LODS_load_string_operand ),
    .o_opcode_x86_LOOP_count ( o_opcode_x86_LOOP_count ),
    .o_opcode_x86_LOOPZ_count_while_zero ( o_opcode_x86_LOOPZ_count_while_zero ),
    .o_opcode_x86_LOOPNZ_count_while_not_zero ( o_opcode_x86_LOOPNZ_count_while_not_zero ),
    .o_opcode_x86_LSL_load_segment_limit ( o_opcode_x86_LSL_load_segment_limit ),
    .o_opcode_x86_LSS_load_pointer_to_SS ( o_opcode_x86_LSS_load_pointer_to_SS ),
    .o_opcode_x86_LTR_load_task_register ( o_opcode_x86_LTR_load_task_register ),
    .o_opcode_x86_MOV_reg_to_reg_mem ( o_opcode_x86_MOV_reg_to_reg_mem ),
    .o_opcode_x86_MOV_reg_mem_to_reg ( o_opcode_x86_MOV_reg_mem_to_reg ),
    .o_opcode_x86_MOV_imm_to_reg_mem ( o_opcode_x86_MOV_imm_to_reg_mem ),
    .o_opcode_x86_MOV_imm_to_reg ( o_opcode_x86_MOV_imm_to_reg ),
    .o_opcode_x86_MOV_mem_to_acc ( o_opcode_x86_MOV_mem_to_acc ),
    .o_opcode_x86_MOV_acc_to_mem ( o_opcode_x86_MOV_acc_to_mem ),
    .o_opcode_x86_MOV_CR_from_reg ( o_opcode_x86_MOV_CR_from_reg ),
    .o_opcode_x86_MOV_reg_from_CR ( o_opcode_x86_MOV_reg_from_CR ),
    .o_opcode_x86_MOV_DR_from_reg ( o_opcode_x86_MOV_DR_from_reg ),
    .o_opcode_x86_MOV_reg_from_DR ( o_opcode_x86_MOV_reg_from_DR ),
    .o_opcode_x86_MOV_TR_from_reg ( o_opcode_x86_MOV_TR_from_reg ),
    .o_opcode_x86_MOV_reg_from_TR ( o_opcode_x86_MOV_reg_from_TR ),
    .o_opcode_x86_MOV_reg_mem_to_sreg ( o_opcode_x86_MOV_reg_mem_to_sreg ),
    .o_opcode_x86_MOV_sreg_to_reg_mem ( o_opcode_x86_MOV_sreg_to_reg_mem ),
    .o_opcode_x86_MOVBE_move_data_after_swapping_bytes_reg_mem_to_reg ( o_opcode_x86_MOVBE_move_data_after_swapping_bytes_reg_mem_to_reg ),
    .o_opcode_x86_MOVBE_move_data_after_swapping_bytes_reg_to_reg_mem ( o_opcode_x86_MOVBE_move_data_after_swapping_bytes_reg_to_reg_mem ),
    .o_opcode_x86_MOVS_move_data_from_string_to_string ( o_opcode_x86_MOVS_move_data_from_string_to_string ),
    .o_opcode_x86_MOVSX_move_with_sign_extend_mem_reg_to_reg ( o_opcode_x86_MOVSX_move_with_sign_extend_mem_reg_to_reg ),
    .o_opcode_x86_MOVZX_move_with_zero_extend_mem_reg_to_reg ( o_opcode_x86_MOVZX_move_with_zero_extend_mem_reg_to_reg ),
    .o_opcode_x86_MUL_acc_with_reg_mem ( o_opcode_x86_MUL_acc_with_reg_mem ),
    .o_opcode_x86_NEG_two_s_complement_negation ( o_opcode_x86_NEG_two_s_complement_negation ),
    .o_opcode_x86_NOP_no_operation ( o_opcode_x86_NOP_no_operation ),
    .o_opcode_x86_NOP_no_operation_multi_byte ( o_opcode_x86_NOP_no_operation_multi_byte ),
    .o_opcode_x86_NOT_one_s_complement_negation ( o_opcode_x86_NOT_one_s_complement_negation ),
    .o_opcode_x86_OR_reg_to_reg_mem ( o_opcode_x86_OR_reg_to_reg_mem ),
    .o_opcode_x86_OR_reg_mem_to_reg ( o_opcode_x86_OR_reg_mem_to_reg ),
    .o_opcode_x86_OR_imm_to_reg_mem ( o_opcode_x86_OR_imm_to_reg_mem ),
    .o_opcode_x86_OR_imm_to_acc ( o_opcode_x86_OR_imm_to_acc ),
    .o_opcode_x86_OUT_port_fixed ( o_opcode_x86_OUT_port_fixed ),
    .o_opcode_x86_OUT_port_variable ( o_opcode_x86_OUT_port_variable ),
    .o_opcode_x86_OUTS_output_string ( o_opcode_x86_OUTS_output_string ),
    .o_opcode_x86_POP_reg_mem ( o_opcode_x86_POP_reg_mem ),
    .o_opcode_x86_POP_reg ( o_opcode_x86_POP_reg ),
    .o_opcode_x86_POP_sreg_2 ( o_opcode_x86_POP_sreg_2 ),
    .o_opcode_x86_POP_sreg_3 ( o_opcode_x86_POP_sreg_3 ),
    .o_opcode_x86_POPA_pop_all_general_registers ( o_opcode_x86_POPA_pop_all_general_registers ),
    .o_opcode_x86_POPF_pop_stack_into_FLAGS_or_EFLAGS ( o_opcode_x86_POPF_pop_stack_into_FLAGS_or_EFLAGS ),
    .o_opcode_x86_PUSH_reg_mem ( o_opcode_x86_PUSH_reg_mem ),
    .o_opcode_x86_PUSH_reg ( o_opcode_x86_PUSH_reg ),
    .o_opcode_x86_PUSH_sreg_2 ( o_opcode_x86_PUSH_sreg_2 ),
    .o_opcode_x86_PUSH_sreg_3 ( o_opcode_x86_PUSH_sreg_3 ),
    .o_opcode_x86_PUSH_imm ( o_opcode_x86_PUSH_imm ),
    .o_opcode_x86_PUSH_all_general_registers ( o_opcode_x86_PUSH_all_general_registers ),
    .o_opcode_x86_PUSHF_push_flags_onto_stack ( o_opcode_x86_PUSHF_push_flags_onto_stack ),
    .o_opcode_x86_RCL_reg_mem_by_1 ( o_opcode_x86_RCL_reg_mem_by_1 ),
    .o_opcode_x86_RCL_reg_mem_by_CL ( o_opcode_x86_RCL_reg_mem_by_CL ),
    .o_opcode_x86_RCL_reg_mem_by_imm ( o_opcode_x86_RCL_reg_mem_by_imm ),
    .o_opcode_x86_RCR_reg_mem_by_1 ( o_opcode_x86_RCR_reg_mem_by_1 ),
    .o_opcode_x86_RCR_reg_mem_by_CL ( o_opcode_x86_RCR_reg_mem_by_CL ),
    .o_opcode_x86_RCR_reg_mem_by_imm ( o_opcode_x86_RCR_reg_mem_by_imm ),
    .o_opcode_x86_RDMSR_read_from_model_specific_reg ( o_opcode_x86_RDMSR_read_from_model_specific_reg ),
    .o_opcode_x86_RDPCM_read_performance_monitoring_counters ( o_opcode_x86_RDPCM_read_performance_monitoring_counters ),
    .o_opcode_x86_RDTSC_read_time_stamp_counter ( o_opcode_x86_RDTSC_read_time_stamp_counter ),
    .o_opcode_x86_RDTSC_read_time_stamp_counter_and_processor_id ( o_opcode_x86_RDTSC_read_time_stamp_counter_and_processor_id ),
    .o_opcode_x86_REP_INS_input_string ( o_opcode_x86_REP_INS_input_string ),
    .o_opcode_x86_REP_LODS_load_string ( o_opcode_x86_REP_LODS_load_string ),
    .o_opcode_x86_REP_MOVS_move_string ( o_opcode_x86_REP_MOVS_move_string ),
    .o_opcode_x86_REP_OUTS_output_string ( o_opcode_x86_REP_OUTS_output_string ),
    .o_opcode_x86_REP_STOS_store_string ( o_opcode_x86_REP_STOS_store_string ),
    .o_opcode_x86_REPE_CMPS_compare_string ( o_opcode_x86_REPE_CMPS_compare_string ),
    .o_opcode_x86_REPE_SCAS_scan_string ( o_opcode_x86_REPE_SCAS_scan_string ),
    .o_opcode_x86_REPNE_CMPS_compare_string ( o_opcode_x86_REPNE_CMPS_compare_string ),
    .o_opcode_x86_REPNE_SCAS_scan_string ( o_opcode_x86_REPNE_SCAS_scan_string ),
    .o_opcode_x86_RET_return_from_procedure_to_same_segment_no_argument ( o_opcode_x86_RET_return_from_procedure_to_same_segment_no_argument ),
    .o_opcode_x86_RET_return_from_procedure_to_same_segment_adding_imm_to_SP ( o_opcode_x86_RET_return_from_procedure_to_same_segment_adding_imm_to_SP ),
    .o_opcode_x86_RET_return_from_procedure_to_other_segment_no_argument ( o_opcode_x86_RET_return_from_procedure_to_other_segment_no_argument ),
    .o_opcode_x86_RET_return_from_procedure_to_other_segment_adding_imm_to_SP ( o_opcode_x86_RET_return_from_procedure_to_other_segment_adding_imm_to_SP ),
    .o_opcode_x86_ROL_reg_mem_by_1 ( o_opcode_x86_ROL_reg_mem_by_1 ),
    .o_opcode_x86_ROL_reg_mem_by_CL ( o_opcode_x86_ROL_reg_mem_by_CL ),
    .o_opcode_x86_ROL_reg_mem_by_imm ( o_opcode_x86_ROL_reg_mem_by_imm ),
    .o_opcode_x86_ROR_reg_mem_by_1 ( o_opcode_x86_ROR_reg_mem_by_1 ),
    .o_opcode_x86_ROR_reg_mem_by_CL ( o_opcode_x86_ROR_reg_mem_by_CL ),
    .o_opcode_x86_ROR_reg_mem_by_imm ( o_opcode_x86_ROR_reg_mem_by_imm ),
    .o_opcode_x86_RSM_resume_from_system_management_mode ( o_opcode_x86_RSM_resume_from_system_management_mode ),
    .o_opcode_x86_SAHF_store_AH_into_flags ( o_opcode_x86_SAHF_store_AH_into_flags ),
    .o_opcode_x86_SAR_reg_mem_by_1 ( o_opcode_x86_SAR_reg_mem_by_1 ),
    .o_opcode_x86_SAR_reg_mem_by_CL ( o_opcode_x86_SAR_reg_mem_by_CL ),
    .o_opcode_x86_SAR_reg_mem_by_imm ( o_opcode_x86_SAR_reg_mem_by_imm ),
    .o_opcode_x86_SBB_reg_to_reg_mem ( o_opcode_x86_SBB_reg_to_reg_mem ),
    .o_opcode_x86_SBB_reg_mem_to_reg ( o_opcode_x86_SBB_reg_mem_to_reg ),
    .o_opcode_x86_SBB_imm_to_reg_mem ( o_opcode_x86_SBB_imm_to_reg_mem ),
    .o_opcode_x86_SBB_imm_to_acc ( o_opcode_x86_SBB_imm_to_acc ),
    .o_opcode_x86_SCAS_scan_string ( o_opcode_x86_SCAS_scan_string ),
    .o_opcode_x86_SETcc_byte_set_on_condition ( o_opcode_x86_SETcc_byte_set_on_condition ),
    .o_opcode_x86_SGDT_store_global_descriptor_table_register ( o_opcode_x86_SGDT_store_global_descriptor_table_register ),
    .o_opcode_x86_SHL_reg_mem_by_1 ( o_opcode_x86_SHL_reg_mem_by_1 ),
    .o_opcode_x86_SHL_reg_mem_by_CL ( o_opcode_x86_SHL_reg_mem_by_CL ),
    .o_opcode_x86_SHL_reg_mem_by_imm ( o_opcode_x86_SHL_reg_mem_by_imm ),
    .o_opcode_x86_SHLD_reg_mem_by_imm ( o_opcode_x86_SHLD_reg_mem_by_imm ),
    .o_opcode_x86_SHLD_reg_mem_by_CL ( o_opcode_x86_SHLD_reg_mem_by_CL ),
    .o_opcode_x86_SHR_reg_mem_by_1 ( o_opcode_x86_SHR_reg_mem_by_1 ),
    .o_opcode_x86_SHR_reg_mem_by_CL ( o_opcode_x86_SHR_reg_mem_by_CL ),
    .o_opcode_x86_SHR_reg_mem_by_imm ( o_opcode_x86_SHR_reg_mem_by_imm ),
    .o_opcode_x86_SHRD_reg_mem_by_imm ( o_opcode_x86_SHRD_reg_mem_by_imm ),
    .o_opcode_x86_SHRD_reg_mem_by_CL ( o_opcode_x86_SHRD_reg_mem_by_CL ),
    .o_opcode_x86_SIDT_store_interrupt_desciptor_table_register ( o_opcode_x86_SIDT_store_interrupt_desciptor_table_register ),
    .o_opcode_x86_SLDT_store_local_desciptor_table_register ( o_opcode_x86_SLDT_store_local_desciptor_table_register ),
    .o_opcode_x86_SMSW_store_machine_status_word ( o_opcode_x86_SMSW_store_machine_status_word ),
    .o_opcode_x86_STC_set_carry_flag ( o_opcode_x86_STC_set_carry_flag ),
    .o_opcode_x86_STD_set_direction_flag ( o_opcode_x86_STD_set_direction_flag ),
    .o_opcode_x86_STI_set_interrupt_enable_flag ( o_opcode_x86_STI_set_interrupt_enable_flag ),
    .o_opcode_x86_STOS_store_string_data ( o_opcode_x86_STOS_store_string_data ),
    .o_opcode_x86_STR_store_task_register ( o_opcode_x86_STR_store_task_register ),
    .o_opcode_x86_SUB_reg_to_reg_mem ( o_opcode_x86_SUB_reg_to_reg_mem ),
    .o_opcode_x86_SUB_reg_mem_to_reg ( o_opcode_x86_SUB_reg_mem_to_reg ),
    .o_opcode_x86_SUB_imm_to_reg_mem ( o_opcode_x86_SUB_imm_to_reg_mem ),
    .o_opcode_x86_SUB_imm_to_acc ( o_opcode_x86_SUB_imm_to_acc ),
    .o_opcode_x86_TEST_reg_mem_and_reg ( o_opcode_x86_TEST_reg_mem_and_reg ),
    .o_opcode_x86_TEST_imm_and_reg_mem ( o_opcode_x86_TEST_imm_and_reg_mem ),
    .o_opcode_x86_TEST_imm_and_acc ( o_opcode_x86_TEST_imm_and_acc ),
    .o_opcode_x86_UD0_undefined_instruction ( o_opcode_x86_UD0_undefined_instruction ),
    .o_opcode_x86_UD1_undefined_instruction ( o_opcode_x86_UD1_undefined_instruction ),
    .o_opcode_x86_UD2_undefined_instruction ( o_opcode_x86_UD2_undefined_instruction ),
    .o_opcode_x86_VERR_verify_a_segment_for_reading ( o_opcode_x86_VERR_verify_a_segment_for_reading ),
    .o_opcode_x86_VERW_verify_a_segment_for_writing ( o_opcode_x86_VERW_verify_a_segment_for_writing ),
    .o_opcode_x86_WAIT_wait ( o_opcode_x86_WAIT_wait ),
    .o_opcode_x86_WBINVD_writeback_and_invalidate_data_cache ( o_opcode_x86_WBINVD_writeback_and_invalidate_data_cache ),
    .o_opcode_x86_WRMSR_write_to_model_specific_register ( o_opcode_x86_WRMSR_write_to_model_specific_register ),
    .o_opcode_x86_XADD_exchange_and_add ( o_opcode_x86_XADD_exchange_and_add ),
    .o_opcode_x86_XCHG_reg_mem_with_reg ( o_opcode_x86_XCHG_reg_mem_with_reg ),
    .o_opcode_x86_XCHG_reg_with_acc_short ( o_opcode_x86_XCHG_reg_with_acc_short ),
    .o_opcode_x86_XLAT_table_look_up_translation ( o_opcode_x86_XLAT_table_look_up_translation ),
    .o_opcode_x86_XOR_reg_to_reg_mem ( o_opcode_x86_XOR_reg_to_reg_mem ),
    .o_opcode_x86_XOR_reg_mem_to_reg ( o_opcode_x86_XOR_reg_mem_to_reg ),
    .o_opcode_x86_XOR_imm_to_reg_mem ( o_opcode_x86_XOR_imm_to_reg_mem ),
    .o_opcode_x86_XOR_imm_to_acc ( o_opcode_x86_XOR_imm_to_acc ),
    .i_instruction ( i_instruction[0:3] )
);

endmodule
