module memory #(
    // parameters
) (
    // port_list
    input  logic [31:0] address,
    input  logic        write_enable,
    input  logic [31:0] write_data,
    input  logic        read_enable,
    output logic [31:0] read_data,
);

// decode_main decode_main_inst (
//     .instruction ( instruction ),
//     .opcode ( opcode ),
//     .operand ( operand ),
// );

endmodule
