/*
project: w80386dx
author: Chang Wei<changwei1006@gmail.com>
repo: https://github.com/openx86/w80386dx
module: decode
create at: 2022-01-04 03:27:51
description: decode module
*/

`include "D:/GitHub/openx86/w80386dx/rtl/definition.h"

module decode (
    output logic        opcode_MOV_reg_to_reg_mem,
    output logic        opcode_MOV_reg_mem_to_reg,
    output logic        opcode_MOV_imm_to_reg_mem,
    output logic        opcode_MOV_imm_to_reg_short,
    output logic        opcode_MOV_mem_to_acc,
    output logic        opcode_MOV_acc_to_mem,
    output logic        opcode_MOV_reg_mem_to_sreg,
    output logic        opcode_MOV_sreg_to_reg_mem,
    output logic        opcode_MOVSX,
    output logic        opcode_MOVZX,
    output logic        opcode_PUSH_reg_mem,
    output logic        opcode_PUSH_reg_short,
    output logic        opcode_PUSH_sreg_2,
    output logic        opcode_PUSH_sreg_3,
    output logic        opcode_PUSH_imm,
    output logic        opcode_PUSH_all,
    output logic        opcode_POP_reg_mem,
    output logic        opcode_POP_reg_short,
    output logic        opcode_POP_sreg_2,
    output logic        opcode_POP_sreg_3,
    output logic        opcode_POP_all,
    output logic        opcode_XCHG_reg_mem_with_reg,
    output logic        opcode_XCHG_reg_with_acc_short,
    output logic        opcode_IN_port_fixed,
    output logic        opcode_IN_port_variable,
    output logic        opcode_OUT_port_fixed,
    output logic        opcode_OUT_port_variable,
    output logic        opcode_LEA_load_ea_to_reg,
    output logic        opcode_LDS_load_ptr_to_DS,
    output logic        opcode_LES_load_ptr_to_ES,
    output logic        opcode_LFS_load_ptr_to_FS,
    output logic        opcode_LGS_load_ptr_to_GS,
    output logic        opcode_LSS_load_ptr_to_SS,
    output logic        opcode_CLC_clear_carry_flag,
    output logic        opcode_CLD_clear_direction_flag,
    output logic        opcode_CLI_clear_interrupt_enable_flag,
    output logic        opcode_CLTS_clear_task_switched_flag,
    output logic        opcode_CMC_complement_carry_flag,
    output logic        opcode_LAHF_load_ah_into_flag,
    output logic        opcode_POPF_pop_flags,
    output logic        opcode_PUSHF_push_flags,
    output logic        opcode_SAHF_store_ah_into_flag,
    output logic        opcode_STC_set_carry_flag,
    output logic        opcode_STD_set_direction_flag,
    output logic        opcode_STI_set_interrupt_enable_flag,
    output logic        opcode_ADD_reg_to_mem,
    output logic        opcode_ADD_mem_to_reg,
    output logic        opcode_ADD_imm_to_reg_mem,
    output logic        opcode_ADD_imm_to_acc,
    output logic        opcode_ADC_reg_to_mem,
    output logic        opcode_ADC_mem_to_reg,
    output logic        opcode_ADC_imm_to_reg_mem,
    output logic        opcode_ADC_imm_to_acc,
    output logic        opcode_INC_reg_mem,
    output logic        opcode_INC_reg,
    output logic        opcode_SUB_reg_to_mem,
    output logic        opcode_SUB_mem_to_reg,
    output logic        opcode_SUB_imm_to_reg_mem,
    output logic        opcode_SUB_imm_to_acc,
    output logic        opcode_SBB_reg_to_mem,
    output logic        opcode_SBB_mem_to_reg,
    output logic        opcode_SBB_imm_to_reg_mem,
    output logic        opcode_SBB_imm_to_acc,
    output logic        opcode_DEC_reg_mem,
    output logic        opcode_DEC_reg,
    output logic        opcode_CMP_mem_with_reg,
    output logic        opcode_CMP_reg_with_mem,
    output logic        opcode_CMP_imm_with_reg_mem,
    output logic        opcode_CMP_imm_with_acc,
    output logic        opcode_NEG_change_sign,
    output logic        opcode_AAA,
    output logic        opcode_AAS,
    output logic        opcode_DAA,
    output logic        opcode_DAS,
    output logic        opcode_MUL_acc_with_reg_mem,
    output logic        opcode_IMUL_acc_with_reg_mem,
    output logic        opcode_IMUL_reg_with_reg_mem,
    output logic        opcode_IMUL_reg_mem_with_imm_to_reg,
    output logic        opcode_DIV_acc_by_reg_mem,
    output logic        opcode_IDIV_acc_by_reg_mem,
    output logic        opcode_AAD,
    output logic        opcode_AAM,
    output logic        opcode_CBW,
    output logic        opcode_CWD,
    output logic        opcode_ROL_reg_mem_by_1,
    output logic        opcode_ROL_reg_mem_by_CL,
    output logic        opcode_ROL_reg_mem_by_imm,
    output logic        opcode_ROR_reg_mem_by_1,
    output logic        opcode_ROR_reg_mem_by_CL,
    output logic        opcode_ROR_reg_mem_by_imm,
    output logic        opcode_SHL_reg_mem_by_1,
    output logic        opcode_SHL_reg_mem_by_CL,
    output logic        opcode_SHL_reg_mem_by_imm,
    output logic        opcode_SAR_reg_mem_by_1,
    output logic        opcode_SAR_reg_mem_by_CL,
    output logic        opcode_SAR_reg_mem_by_imm,
    output logic        opcode_SHR_reg_mem_by_1,
    output logic        opcode_SHR_reg_mem_by_CL,
    output logic        opcode_SHR_reg_mem_by_imm,
    output logic        opcode_RCL_reg_mem_by_1,
    output logic        opcode_RCL_reg_mem_by_CL,
    output logic        opcode_RCL_reg_mem_by_imm,
    output logic        opcode_RCR_reg_mem_by_1,
    output logic        opcode_RCR_reg_mem_by_CL,
    output logic        opcode_RCR_reg_mem_by_imm,
    output logic        opcode_SHLD_reg_mem_by_imm,
    output logic        opcode_SHLD_reg_mem_by_CL,
    output logic        opcode_SHRD_reg_mem_by_imm,
    output logic        opcode_SHRD_reg_mem_by_CL,
    output logic        opcode_AND_reg_to_mem,
    output logic        opcode_AND_mem_to_reg,
    output logic        opcode_AND_imm_to_reg_mem,
    output logic        opcode_AND_imm_to_acc,
    output logic        opcode_TEST_reg_mem_and_reg,
    output logic        opcode_TEST_imm_to_reg_mem,
    output logic        opcode_TEST_imm_to_acc,
    output logic        opcode_OR_reg_to_mem,
    output logic        opcode_OR_mem_to_reg,
    output logic        opcode_OR_imm_to_reg_mem,
    output logic        opcode_OR_imm_to_acc,
    output logic        opcode_XOR_reg_to_mem,
    output logic        opcode_XOR_mem_to_reg,
    output logic        opcode_XOR_imm_to_reg_mem,
    output logic        opcode_XOR_imm_to_acc,
    output logic        opcode_NOT,
    output logic        opcode_CMPS,
    output logic        opcode_INS,
    output logic        opcode_LODS,
    output logic        opcode_MOVS,
    output logic        opcode_OUTS,
    output logic        opcode_SCAS,
    output logic        opcode_STOS,
    output logic        opcode_XLAT,
    output logic        opcode_REPE,
    output logic        opcode_REPNE,
    output logic        opcode_BSF,
    output logic        opcode_BSR,
    output logic        opcode_BT_reg_mem_with_imm,
    output logic        opcode_BT_reg_mem_with_reg,
    output logic        opcode_BTC_reg_mem_with_imm,
    output logic        opcode_BTC_reg_mem_with_reg,
    output logic        opcode_BTR_reg_mem_with_imm,
    output logic        opcode_BTR_reg_mem_with_reg,
    output logic        opcode_BTS_reg_mem_with_imm,
    output logic        opcode_BTS_reg_mem_with_reg,
    output logic        opcode_CALL_direct_within_segment,
    output logic        opcode_CALL_indirect_within_segment,
    output logic        opcode_CALL_direct_intersegment,
    output logic        opcode_CALL_indirect_intersegment,
    output logic        opcode_JMP_short,
    output logic        opcode_JMP_direct_within_segment,
    output logic        opcode_JMP_indirect_within_segment,
    output logic        opcode_JMP_direct_intersegment,
    output logic        opcode_JMP_indirect_intersegment,
    output logic        opcode_RET_within_segment,
    output logic        opcode_RET_within_segment_adding_imm_to_SP,
    output logic        opcode_RET_intersegment,
    output logic        opcode_RET_intersegment_adding_imm_to_SP,
    output logic        opcode_JO_8bit_disp,
    output logic        opcode_JO_full_disp,
    output logic        opcode_JNO_8bit_disp,
    output logic        opcode_JNO_full_disp,
    output logic        opcode_JB_8bit_disp,
    output logic        opcode_JB_full_disp,
    output logic        opcode_JNB_8bit_disp,
    output logic        opcode_JNB_full_disp,
    output logic        opcode_JE_8bit_disp,
    output logic        opcode_JE_full_disp,
    output logic        opcode_JNE_8bit_disp,
    output logic        opcode_JNE_full_disp,
    output logic        opcode_JBE_8bit_disp,
    output logic        opcode_JBE_full_disp,
    output logic        opcode_JNBE_8bit_disp,
    output logic        opcode_JNBE_full_disp,
    output logic        opcode_JS_8bit_disp,
    output logic        opcode_JS_full_disp,
    output logic        opcode_JNS_8bit_disp,
    output logic        opcode_JNS_full_disp,
    output logic        opcode_JP_8bit_disp,
    output logic        opcode_JP_full_disp,
    output logic        opcode_JNP_8bit_disp,
    output logic        opcode_JNP_full_disp,
    output logic        opcode_JL_8bit_disp,
    output logic        opcode_JL_full_disp,
    output logic        opcode_JNL_8bit_disp,
    output logic        opcode_JNL_full_disp,
    output logic        opcode_JLE_8bit_disp,
    output logic        opcode_JLE_full_disp,
    output logic        opcode_JNLE_8bit_disp,
    output logic        opcode_JNLE_full_disp,
    output logic        opcode_JCXZ,
    output logic        opcode_LOOP,
    output logic        opcode_LOOPZ,
    output logic        opcode_LOOPNZ,
    output logic        opcode_SETO,
    output logic        opcode_SETNO,
    output logic        opcode_SETB,
    output logic        opcode_SETNB,
    output logic        opcode_SETE,
    output logic        opcode_SETNE,
    output logic        opcode_SETBE,
    output logic        opcode_SETNBE,
    output logic        opcode_SETS,
    output logic        opcode_SETNS,
    output logic        opcode_SETP,
    output logic        opcode_SETNP,
    output logic        opcode_SETL,
    output logic        opcode_SETNL,
    output logic        opcode_SETLE,
    output logic        opcode_SETNLE,
    output logic        opcode_ENTER,
    output logic        opcode_LEAVE,
    output logic        opcode_INT_type_3,
    output logic        opcode_INT_type_specified,
    output logic        opcode_INTO,
    output logic        opcode_BOUND,
    output logic        opcode_IRET,
    output logic        opcode_HLT,
    output logic        opcode_MOV_CR0_CR2_CR3_from_reg,
    output logic        opcode_MOV_reg_from_CR0_3,
    output logic        opcode_MOV_DR0_7_from_reg,
    output logic        opcode_MOV_reg_from_DR0_7,
    output logic        opcode_MOV_TR6_7_from_reg,
    output logic        opcode_MOV_reg_from_TR6_7,
    output logic        opcode_NOP,
    output logic        opcode_WAIT,
    output logic        opcode_processor_extension_escape,
    output logic        opcode_prefix_address_size,
    output logic        opcode_prefix_bus_lock,
    output logic        opcode_prefix_operand_size,
    output logic        opcode_prefix_segment_override_CS,
    output logic        opcode_prefix_segment_override_DS,
    output logic        opcode_prefix_segment_override_ES,
    output logic        opcode_prefix_segment_override_FS,
    output logic        opcode_prefix_segment_override_GS,
    output logic        opcode_prefix_segment_override_SS,
    output logic        opcode_ARPL,
    output logic        opcode_LAR,
    output logic        opcode_LGDT,
    output logic        opcode_LIDT,
    output logic        opcode_LLDT,
    output logic        opcode_LMSW,
    output logic        opcode_LSL,
    output logic        opcode_LTR,
    output logic        opcode_SGDT,
    output logic        opcode_SIDT,
    output logic        opcode_SLDT,
    output logic        opcode_SMSW,
    output logic        opcode_STR,
    output logic        opcode_VERR,
    output logic        opcode_VERW,
    // input  logic [`info_bit_width_len-1:0] bit_width,
    // output logic [`info_reg_seg_len-1:0] info_segment_reg,
    // output logic [`info_reg_gpr_len-1:0] info_base_reg,
    // output logic [`info_reg_gpr_len-1:0] info_index_reg,
    // output logic [`info_displacement_len-1:0] info_displacement,
    // output logic        sib_is_present,
    // output logic [ 3:0] instruction_length,
    input  logic [ 7:0] instruction [0:9]
);

// logic        s;
// logic        w;
// logic [ 2:0] gereral_propose_register;
// logic [ 2:0] sreg;
// logic [ 1:0] mod;
// logic [ 2:0] rm;
// logic        has_s;
// logic        has_w;
// logic        has_sreg;
// logic        has_mod_rm;
// logic        is_prefix_segment;
// logic        is_prefix;

decode_opcode u_decode_opcode (
    .opcode_MOV_reg_to_reg_mem ( opcode_MOV_reg_to_reg_mem ),
    .opcode_MOV_reg_mem_to_reg ( opcode_MOV_reg_mem_to_reg ),
    .opcode_MOV_imm_to_reg_mem ( opcode_MOV_imm_to_reg_mem ),
    .opcode_MOV_imm_to_reg_short ( opcode_MOV_imm_to_reg_short ),
    .opcode_MOV_mem_to_acc ( opcode_MOV_mem_to_acc ),
    .opcode_MOV_acc_to_mem ( opcode_MOV_acc_to_mem ),
    .opcode_MOV_reg_mem_to_sreg ( opcode_MOV_reg_mem_to_sreg ),
    .opcode_MOV_sreg_to_reg_mem ( opcode_MOV_sreg_to_reg_mem ),
    .opcode_MOVSX ( opcode_MOVSX ),
    .opcode_MOVZX ( opcode_MOVZX ),
    .opcode_PUSH_reg_mem ( opcode_PUSH_reg_mem ),
    .opcode_PUSH_reg_short ( opcode_PUSH_reg_short ),
    .opcode_PUSH_sreg_2 ( opcode_PUSH_sreg_2 ),
    .opcode_PUSH_sreg_3 ( opcode_PUSH_sreg_3 ),
    .opcode_PUSH_imm ( opcode_PUSH_imm ),
    .opcode_PUSH_all ( opcode_PUSH_all ),
    .opcode_POP_reg_mem ( opcode_POP_reg_mem ),
    .opcode_POP_reg_short ( opcode_POP_reg_short ),
    .opcode_POP_sreg_2 ( opcode_POP_sreg_2 ),
    .opcode_POP_sreg_3 ( opcode_POP_sreg_3 ),
    .opcode_POP_all ( opcode_POP_all ),
    .opcode_XCHG_reg_mem_with_reg ( opcode_XCHG_reg_mem_with_reg ),
    .opcode_XCHG_reg_with_acc_short ( opcode_XCHG_reg_with_acc_short ),
    .opcode_IN_port_fixed ( opcode_IN_port_fixed ),
    .opcode_IN_port_variable ( opcode_IN_port_variable ),
    .opcode_OUT_port_fixed ( opcode_OUT_port_fixed ),
    .opcode_OUT_port_variable ( opcode_OUT_port_variable ),
    .opcode_LEA_load_ea_to_reg ( opcode_LEA_load_ea_to_reg ),
    .opcode_LDS_load_ptr_to_DS ( opcode_LDS_load_ptr_to_DS ),
    .opcode_LES_load_ptr_to_ES ( opcode_LES_load_ptr_to_ES ),
    .opcode_LFS_load_ptr_to_FS ( opcode_LFS_load_ptr_to_FS ),
    .opcode_LGS_load_ptr_to_GS ( opcode_LGS_load_ptr_to_GS ),
    .opcode_LSS_load_ptr_to_SS ( opcode_LSS_load_ptr_to_SS ),
    .opcode_CLC_clear_carry_flag ( opcode_CLC_clear_carry_flag ),
    .opcode_CLD_clear_direction_flag ( opcode_CLD_clear_direction_flag ),
    .opcode_CLI_clear_interrupt_enable_flag ( opcode_CLI_clear_interrupt_enable_flag ),
    .opcode_CLTS_clear_task_switched_flag ( opcode_CLTS_clear_task_switched_flag ),
    .opcode_CMC_complement_carry_flag ( opcode_CMC_complement_carry_flag ),
    .opcode_LAHF_load_ah_into_flag ( opcode_LAHF_load_ah_into_flag ),
    .opcode_POPF_pop_flags ( opcode_POPF_pop_flags ),
    .opcode_PUSHF_push_flags ( opcode_PUSHF_push_flags ),
    .opcode_SAHF_store_ah_into_flag ( opcode_SAHF_store_ah_into_flag ),
    .opcode_STC_set_carry_flag ( opcode_STC_set_carry_flag ),
    .opcode_STD_set_direction_flag ( opcode_STD_set_direction_flag ),
    .opcode_STI_set_interrupt_enable_flag ( opcode_STI_set_interrupt_enable_flag ),
    .opcode_ADD_reg_to_mem ( opcode_ADD_reg_to_mem ),
    .opcode_ADD_mem_to_reg ( opcode_ADD_mem_to_reg ),
    .opcode_ADD_imm_to_reg_mem ( opcode_ADD_imm_to_reg_mem ),
    .opcode_ADD_imm_to_acc ( opcode_ADD_imm_to_acc ),
    .opcode_ADC_reg_to_mem ( opcode_ADC_reg_to_mem ),
    .opcode_ADC_mem_to_reg ( opcode_ADC_mem_to_reg ),
    .opcode_ADC_imm_to_reg_mem ( opcode_ADC_imm_to_reg_mem ),
    .opcode_ADC_imm_to_acc ( opcode_ADC_imm_to_acc ),
    .opcode_INC_reg_mem ( opcode_INC_reg_mem ),
    .opcode_INC_reg ( opcode_INC_reg ),
    .opcode_SUB_reg_to_mem ( opcode_SUB_reg_to_mem ),
    .opcode_SUB_mem_to_reg ( opcode_SUB_mem_to_reg ),
    .opcode_SUB_imm_to_reg_mem ( opcode_SUB_imm_to_reg_mem ),
    .opcode_SUB_imm_to_acc ( opcode_SUB_imm_to_acc ),
    .opcode_SBB_reg_to_mem ( opcode_SBB_reg_to_mem ),
    .opcode_SBB_mem_to_reg ( opcode_SBB_mem_to_reg ),
    .opcode_SBB_imm_to_reg_mem ( opcode_SBB_imm_to_reg_mem ),
    .opcode_SBB_imm_to_acc ( opcode_SBB_imm_to_acc ),
    .opcode_DEC_reg_mem ( opcode_DEC_reg_mem ),
    .opcode_DEC_reg ( opcode_DEC_reg ),
    .opcode_CMP_mem_with_reg ( opcode_CMP_mem_with_reg ),
    .opcode_CMP_reg_with_mem ( opcode_CMP_reg_with_mem ),
    .opcode_CMP_imm_with_reg_mem ( opcode_CMP_imm_with_reg_mem ),
    .opcode_CMP_imm_with_acc ( opcode_CMP_imm_with_acc ),
    .opcode_NEG_change_sign ( opcode_NEG_change_sign ),
    .opcode_AAA ( opcode_AAA ),
    .opcode_AAS ( opcode_AAS ),
    .opcode_DAA ( opcode_DAA ),
    .opcode_DAS ( opcode_DAS ),
    .opcode_MUL_acc_with_reg_mem ( opcode_MUL_acc_with_reg_mem ),
    .opcode_IMUL_acc_with_reg_mem ( opcode_IMUL_acc_with_reg_mem ),
    .opcode_IMUL_reg_with_reg_mem ( opcode_IMUL_reg_with_reg_mem ),
    .opcode_IMUL_reg_mem_with_imm_to_reg ( opcode_IMUL_reg_mem_with_imm_to_reg ),
    .opcode_DIV_acc_by_reg_mem ( opcode_DIV_acc_by_reg_mem ),
    .opcode_IDIV_acc_by_reg_mem ( opcode_IDIV_acc_by_reg_mem ),
    .opcode_AAD ( opcode_AAD ),
    .opcode_AAM ( opcode_AAM ),
    .opcode_CBW ( opcode_CBW ),
    .opcode_CWD ( opcode_CWD ),
    .opcode_ROL_reg_mem_by_1 ( opcode_ROL_reg_mem_by_1 ),
    .opcode_ROL_reg_mem_by_CL ( opcode_ROL_reg_mem_by_CL ),
    .opcode_ROL_reg_mem_by_imm ( opcode_ROL_reg_mem_by_imm ),
    .opcode_ROR_reg_mem_by_1 ( opcode_ROR_reg_mem_by_1 ),
    .opcode_ROR_reg_mem_by_CL ( opcode_ROR_reg_mem_by_CL ),
    .opcode_ROR_reg_mem_by_imm ( opcode_ROR_reg_mem_by_imm ),
    .opcode_SHL_reg_mem_by_1 ( opcode_SHL_reg_mem_by_1 ),
    .opcode_SHL_reg_mem_by_CL ( opcode_SHL_reg_mem_by_CL ),
    .opcode_SHL_reg_mem_by_imm ( opcode_SHL_reg_mem_by_imm ),
    .opcode_SAR_reg_mem_by_1 ( opcode_SAR_reg_mem_by_1 ),
    .opcode_SAR_reg_mem_by_CL ( opcode_SAR_reg_mem_by_CL ),
    .opcode_SAR_reg_mem_by_imm ( opcode_SAR_reg_mem_by_imm ),
    .opcode_SHR_reg_mem_by_1 ( opcode_SHR_reg_mem_by_1 ),
    .opcode_SHR_reg_mem_by_CL ( opcode_SHR_reg_mem_by_CL ),
    .opcode_SHR_reg_mem_by_imm ( opcode_SHR_reg_mem_by_imm ),
    .opcode_RCL_reg_mem_by_1 ( opcode_RCL_reg_mem_by_1 ),
    .opcode_RCL_reg_mem_by_CL ( opcode_RCL_reg_mem_by_CL ),
    .opcode_RCL_reg_mem_by_imm ( opcode_RCL_reg_mem_by_imm ),
    .opcode_RCR_reg_mem_by_1 ( opcode_RCR_reg_mem_by_1 ),
    .opcode_RCR_reg_mem_by_CL ( opcode_RCR_reg_mem_by_CL ),
    .opcode_RCR_reg_mem_by_imm ( opcode_RCR_reg_mem_by_imm ),
    .opcode_SHLD_reg_mem_by_imm ( opcode_SHLD_reg_mem_by_imm ),
    .opcode_SHLD_reg_mem_by_CL ( opcode_SHLD_reg_mem_by_CL ),
    .opcode_SHRD_reg_mem_by_imm ( opcode_SHRD_reg_mem_by_imm ),
    .opcode_SHRD_reg_mem_by_CL ( opcode_SHRD_reg_mem_by_CL ),
    .opcode_AND_reg_to_mem ( opcode_AND_reg_to_mem ),
    .opcode_AND_mem_to_reg ( opcode_AND_mem_to_reg ),
    .opcode_AND_imm_to_reg_mem ( opcode_AND_imm_to_reg_mem ),
    .opcode_AND_imm_to_acc ( opcode_AND_imm_to_acc ),
    .opcode_TEST_reg_mem_and_reg ( opcode_TEST_reg_mem_and_reg ),
    .opcode_TEST_imm_to_reg_mem ( opcode_TEST_imm_to_reg_mem ),
    .opcode_TEST_imm_to_acc ( opcode_TEST_imm_to_acc ),
    .opcode_OR_reg_to_mem ( opcode_OR_reg_to_mem ),
    .opcode_OR_mem_to_reg ( opcode_OR_mem_to_reg ),
    .opcode_OR_imm_to_reg_mem ( opcode_OR_imm_to_reg_mem ),
    .opcode_OR_imm_to_acc ( opcode_OR_imm_to_acc ),
    .opcode_XOR_reg_to_mem ( opcode_XOR_reg_to_mem ),
    .opcode_XOR_mem_to_reg ( opcode_XOR_mem_to_reg ),
    .opcode_XOR_imm_to_reg_mem ( opcode_XOR_imm_to_reg_mem ),
    .opcode_XOR_imm_to_acc ( opcode_XOR_imm_to_acc ),
    .opcode_NOT ( opcode_NOT ),
    .opcode_CMPS ( opcode_CMPS ),
    .opcode_INS ( opcode_INS ),
    .opcode_LODS ( opcode_LODS ),
    .opcode_MOVS ( opcode_MOVS ),
    .opcode_OUTS ( opcode_OUTS ),
    .opcode_SCAS ( opcode_SCAS ),
    .opcode_STOS ( opcode_STOS ),
    .opcode_XLAT ( opcode_XLAT ),
    .opcode_REPE ( opcode_REPE ),
    .opcode_REPNE ( opcode_REPNE ),
    .opcode_BSF ( opcode_BSF ),
    .opcode_BSR ( opcode_BSR ),
    .opcode_BT_reg_mem_with_imm ( opcode_BT_reg_mem_with_imm ),
    .opcode_BT_reg_mem_with_reg ( opcode_BT_reg_mem_with_reg ),
    .opcode_BTC_reg_mem_with_imm ( opcode_BTC_reg_mem_with_imm ),
    .opcode_BTC_reg_mem_with_reg ( opcode_BTC_reg_mem_with_reg ),
    .opcode_BTR_reg_mem_with_imm ( opcode_BTR_reg_mem_with_imm ),
    .opcode_BTR_reg_mem_with_reg ( opcode_BTR_reg_mem_with_reg ),
    .opcode_BTS_reg_mem_with_imm ( opcode_BTS_reg_mem_with_imm ),
    .opcode_BTS_reg_mem_with_reg ( opcode_BTS_reg_mem_with_reg ),
    .opcode_CALL_direct_within_segment ( opcode_CALL_direct_within_segment ),
    .opcode_CALL_indirect_within_segment ( opcode_CALL_indirect_within_segment ),
    .opcode_CALL_direct_intersegment ( opcode_CALL_direct_intersegment ),
    .opcode_CALL_indirect_intersegment ( opcode_CALL_indirect_intersegment ),
    .opcode_JMP_short ( opcode_JMP_short ),
    .opcode_JMP_direct_within_segment ( opcode_JMP_direct_within_segment ),
    .opcode_JMP_indirect_within_segment ( opcode_JMP_indirect_within_segment ),
    .opcode_JMP_direct_intersegment ( opcode_JMP_direct_intersegment ),
    .opcode_JMP_indirect_intersegment ( opcode_JMP_indirect_intersegment ),
    .opcode_RET_within_segment ( opcode_RET_within_segment ),
    .opcode_RET_within_segment_adding_imm_to_SP ( opcode_RET_within_segment_adding_imm_to_SP ),
    .opcode_RET_intersegment ( opcode_RET_intersegment ),
    .opcode_RET_intersegment_adding_imm_to_SP ( opcode_RET_intersegment_adding_imm_to_SP ),
    .opcode_JO_8bit_disp ( opcode_JO_8bit_disp ),
    .opcode_JO_full_disp ( opcode_JO_full_disp ),
    .opcode_JNO_8bit_disp ( opcode_JNO_8bit_disp ),
    .opcode_JNO_full_disp ( opcode_JNO_full_disp ),
    .opcode_JB_8bit_disp ( opcode_JB_8bit_disp ),
    .opcode_JB_full_disp ( opcode_JB_full_disp ),
    .opcode_JNB_8bit_disp ( opcode_JNB_8bit_disp ),
    .opcode_JNB_full_disp ( opcode_JNB_full_disp ),
    .opcode_JE_8bit_disp ( opcode_JE_8bit_disp ),
    .opcode_JE_full_disp ( opcode_JE_full_disp ),
    .opcode_JNE_8bit_disp ( opcode_JNE_8bit_disp ),
    .opcode_JNE_full_disp ( opcode_JNE_full_disp ),
    .opcode_JBE_8bit_disp ( opcode_JBE_8bit_disp ),
    .opcode_JBE_full_disp ( opcode_JBE_full_disp ),
    .opcode_JNBE_8bit_disp ( opcode_JNBE_8bit_disp ),
    .opcode_JNBE_full_disp ( opcode_JNBE_full_disp ),
    .opcode_JS_8bit_disp ( opcode_JS_8bit_disp ),
    .opcode_JS_full_disp ( opcode_JS_full_disp ),
    .opcode_JNS_8bit_disp ( opcode_JNS_8bit_disp ),
    .opcode_JNS_full_disp ( opcode_JNS_full_disp ),
    .opcode_JP_8bit_disp ( opcode_JP_8bit_disp ),
    .opcode_JP_full_disp ( opcode_JP_full_disp ),
    .opcode_JNP_8bit_disp ( opcode_JNP_8bit_disp ),
    .opcode_JNP_full_disp ( opcode_JNP_full_disp ),
    .opcode_JL_8bit_disp ( opcode_JL_8bit_disp ),
    .opcode_JL_full_disp ( opcode_JL_full_disp ),
    .opcode_JNL_8bit_disp ( opcode_JNL_8bit_disp ),
    .opcode_JNL_full_disp ( opcode_JNL_full_disp ),
    .opcode_JLE_8bit_disp ( opcode_JLE_8bit_disp ),
    .opcode_JLE_full_disp ( opcode_JLE_full_disp ),
    .opcode_JNLE_8bit_disp ( opcode_JNLE_8bit_disp ),
    .opcode_JNLE_full_disp ( opcode_JNLE_full_disp ),
    .opcode_JCXZ ( opcode_JCXZ ),
    .opcode_LOOP ( opcode_LOOP ),
    .opcode_LOOPZ ( opcode_LOOPZ ),
    .opcode_LOOPNZ ( opcode_LOOPNZ ),
    .opcode_SETO ( opcode_SETO ),
    .opcode_SETNO ( opcode_SETNO ),
    .opcode_SETB ( opcode_SETB ),
    .opcode_SETNB ( opcode_SETNB ),
    .opcode_SETE ( opcode_SETE ),
    .opcode_SETNE ( opcode_SETNE ),
    .opcode_SETBE ( opcode_SETBE ),
    .opcode_SETNBE ( opcode_SETNBE ),
    .opcode_SETS ( opcode_SETS ),
    .opcode_SETNS ( opcode_SETNS ),
    .opcode_SETP ( opcode_SETP ),
    .opcode_SETNP ( opcode_SETNP ),
    .opcode_SETL ( opcode_SETL ),
    .opcode_SETNL ( opcode_SETNL ),
    .opcode_SETLE ( opcode_SETLE ),
    .opcode_SETNLE ( opcode_SETNLE ),
    .opcode_ENTER ( opcode_ENTER ),
    .opcode_LEAVE ( opcode_LEAVE ),
    .opcode_INT_type_3 ( opcode_INT_type_3 ),
    .opcode_INT_type_specified ( opcode_INT_type_specified ),
    .opcode_INTO ( opcode_INTO ),
    .opcode_BOUND ( opcode_BOUND ),
    .opcode_IRET ( opcode_IRET ),
    .opcode_HLT ( opcode_HLT ),
    .opcode_MOV_CR0_CR2_CR3_from_reg ( opcode_MOV_CR0_CR2_CR3_from_reg ),
    .opcode_MOV_reg_from_CR0_3 ( opcode_MOV_reg_from_CR0_3 ),
    .opcode_MOV_DR0_7_from_reg ( opcode_MOV_DR0_7_from_reg ),
    .opcode_MOV_reg_from_DR0_7 ( opcode_MOV_reg_from_DR0_7 ),
    .opcode_MOV_TR6_7_from_reg ( opcode_MOV_TR6_7_from_reg ),
    .opcode_MOV_reg_from_TR6_7 ( opcode_MOV_reg_from_TR6_7 ),
    .opcode_NOP ( opcode_NOP ),
    .opcode_WAIT ( opcode_WAIT ),
    .opcode_processor_extension_escape ( opcode_processor_extension_escape ),
    .opcode_prefix_address_size ( opcode_prefix_address_size ),
    .opcode_prefix_bus_lock ( opcode_prefix_bus_lock ),
    .opcode_prefix_operand_size ( opcode_prefix_operand_size ),
    .opcode_prefix_segment_override_CS ( opcode_prefix_segment_override_CS ),
    .opcode_prefix_segment_override_DS ( opcode_prefix_segment_override_DS ),
    .opcode_prefix_segment_override_ES ( opcode_prefix_segment_override_ES ),
    .opcode_prefix_segment_override_FS ( opcode_prefix_segment_override_FS ),
    .opcode_prefix_segment_override_GS ( opcode_prefix_segment_override_GS ),
    .opcode_prefix_segment_override_SS ( opcode_prefix_segment_override_SS ),
    .opcode_ARPL ( opcode_ARPL ),
    .opcode_LAR ( opcode_LAR ),
    .opcode_LGDT ( opcode_LGDT ),
    .opcode_LIDT ( opcode_LIDT ),
    .opcode_LLDT ( opcode_LLDT ),
    .opcode_LMSW ( opcode_LMSW ),
    .opcode_LSL ( opcode_LSL ),
    .opcode_LTR ( opcode_LTR ),
    .opcode_SGDT ( opcode_SGDT ),
    .opcode_SIDT ( opcode_SIDT ),
    .opcode_SLDT ( opcode_SLDT ),
    .opcode_SMSW ( opcode_SMSW ),
    .opcode_STR ( opcode_STR ),
    .opcode_VERR ( opcode_VERR ),
    .opcode_VERW ( opcode_VERW ),
    .instruction ( instruction[0:2] )
);

// decode_field u_decode_field (
//     .opcode_MOV_reg_to_reg_mem ( opcode_MOV_reg_to_reg_mem ),
//     .opcode_MOV_reg_mem_to_reg ( opcode_MOV_reg_mem_to_reg ),
//     .opcode_MOV_imm_to_reg_mem ( opcode_MOV_imm_to_reg_mem ),
//     .opcode_MOV_imm_to_reg_short ( opcode_MOV_imm_to_reg_short ),
//     .opcode_MOV_mem_to_acc ( opcode_MOV_mem_to_acc ),
//     .opcode_MOV_acc_to_mem ( opcode_MOV_acc_to_mem ),
//     .opcode_MOV_reg_mem_to_sreg ( opcode_MOV_reg_mem_to_sreg ),
//     .opcode_MOV_sreg_to_reg_mem ( opcode_MOV_sreg_to_reg_mem ),
//     .opcode_MOVSX ( opcode_MOVSX ),
//     .opcode_MOVZX ( opcode_MOVZX ),
//     .opcode_PUSH_reg_mem ( opcode_PUSH_reg_mem ),
//     .opcode_PUSH_reg_short ( opcode_PUSH_reg_short ),
//     .opcode_PUSH_sreg_2 ( opcode_PUSH_sreg_2 ),
//     .opcode_PUSH_sreg_3 ( opcode_PUSH_sreg_3 ),
//     .opcode_PUSH_imm ( opcode_PUSH_imm ),
//     .opcode_PUSH_all ( opcode_PUSH_all ),
//     .opcode_POP_reg_mem ( opcode_POP_reg_mem ),
//     .opcode_POP_reg_short ( opcode_POP_reg_short ),
//     .opcode_POP_sreg_2 ( opcode_POP_sreg_2 ),
//     .opcode_POP_sreg_3 ( opcode_POP_sreg_3 ),
//     .opcode_POP_all ( opcode_POP_all ),
//     .opcode_XCHG_reg_mem_with_reg ( opcode_XCHG_reg_mem_with_reg ),
//     .opcode_XCHG_reg_with_acc_short ( opcode_XCHG_reg_with_acc_short ),
//     .opcode_IN_port_fixed ( opcode_IN_port_fixed ),
//     .opcode_IN_port_variable ( opcode_IN_port_variable ),
//     .opcode_OUT_port_fixed ( opcode_OUT_port_fixed ),
//     .opcode_OUT_port_variable ( opcode_OUT_port_variable ),
//     .opcode_LEA_load_ea_to_reg ( opcode_LEA_load_ea_to_reg ),
//     .opcode_LDS_load_ptr_to_DS ( opcode_LDS_load_ptr_to_DS ),
//     .opcode_LES_load_ptr_to_ES ( opcode_LES_load_ptr_to_ES ),
//     .opcode_LFS_load_ptr_to_FS ( opcode_LFS_load_ptr_to_FS ),
//     .opcode_LGS_load_ptr_to_GS ( opcode_LGS_load_ptr_to_GS ),
//     .opcode_LSS_load_ptr_to_SS ( opcode_LSS_load_ptr_to_SS ),
//     .opcode_CLC_clear_carry_flag ( opcode_CLC_clear_carry_flag ),
//     .opcode_CLD_clear_direction_flag ( opcode_CLD_clear_direction_flag ),
//     .opcode_CLI_clear_interrupt_enable_flag ( opcode_CLI_clear_interrupt_enable_flag ),
//     .opcode_CLTS_clear_task_switched_flag ( opcode_CLTS_clear_task_switched_flag ),
//     .opcode_CMC_complement_carry_flag ( opcode_CMC_complement_carry_flag ),
//     .opcode_LAHF_load_ah_into_flag ( opcode_LAHF_load_ah_into_flag ),
//     .opcode_POPF_pop_flags ( opcode_POPF_pop_flags ),
//     .opcode_PUSHF_push_flags ( opcode_PUSHF_push_flags ),
//     .opcode_SAHF_store_ah_into_flag ( opcode_SAHF_store_ah_into_flag ),
//     .opcode_STC_set_carry_flag ( opcode_STC_set_carry_flag ),
//     .opcode_STD_set_direction_flag ( opcode_STD_set_direction_flag ),
//     .opcode_STI_set_interrupt_enable_flag ( opcode_STI_set_interrupt_enable_flag ),
//     .opcode_ADD_reg_to_mem ( opcode_ADD_reg_to_mem ),
//     .opcode_ADD_mem_to_reg ( opcode_ADD_mem_to_reg ),
//     .opcode_ADD_imm_to_reg_mem ( opcode_ADD_imm_to_reg_mem ),
//     .opcode_ADD_imm_to_acc ( opcode_ADD_imm_to_acc ),
//     .opcode_ADC_reg_to_mem ( opcode_ADC_reg_to_mem ),
//     .opcode_ADC_mem_to_reg ( opcode_ADC_mem_to_reg ),
//     .opcode_ADC_imm_to_reg_mem ( opcode_ADC_imm_to_reg_mem ),
//     .opcode_ADC_imm_to_acc ( opcode_ADC_imm_to_acc ),
//     .opcode_INC_reg_mem ( opcode_INC_reg_mem ),
//     .opcode_INC_reg ( opcode_INC_reg ),
//     .opcode_SUB_reg_to_mem ( opcode_SUB_reg_to_mem ),
//     .opcode_SUB_mem_to_reg ( opcode_SUB_mem_to_reg ),
//     .opcode_SUB_imm_to_reg_mem ( opcode_SUB_imm_to_reg_mem ),
//     .opcode_SUB_imm_to_acc ( opcode_SUB_imm_to_acc ),
//     .opcode_SBB_reg_to_mem ( opcode_SBB_reg_to_mem ),
//     .opcode_SBB_mem_to_reg ( opcode_SBB_mem_to_reg ),
//     .opcode_SBB_imm_to_reg_mem ( opcode_SBB_imm_to_reg_mem ),
//     .opcode_SBB_imm_to_acc ( opcode_SBB_imm_to_acc ),
//     .opcode_DEC_reg_mem ( opcode_DEC_reg_mem ),
//     .opcode_DEC_reg ( opcode_DEC_reg ),
//     .opcode_CMP_mem_with_reg ( opcode_CMP_mem_with_reg ),
//     .opcode_CMP_reg_with_mem ( opcode_CMP_reg_with_mem ),
//     .opcode_CMP_imm_with_reg_mem ( opcode_CMP_imm_with_reg_mem ),
//     .opcode_CMP_imm_with_acc ( opcode_CMP_imm_with_acc ),
//     .opcode_NEG_change_sign ( opcode_NEG_change_sign ),
//     .opcode_AAA ( opcode_AAA ),
//     .opcode_AAS ( opcode_AAS ),
//     .opcode_DAA ( opcode_DAA ),
//     .opcode_DAS ( opcode_DAS ),
//     .opcode_MUL_acc_with_reg_mem ( opcode_MUL_acc_with_reg_mem ),
//     .opcode_IMUL_acc_with_reg_mem ( opcode_IMUL_acc_with_reg_mem ),
//     .opcode_IMUL_reg_with_reg_mem ( opcode_IMUL_reg_with_reg_mem ),
//     .opcode_IMUL_reg_mem_with_imm_to_reg ( opcode_IMUL_reg_mem_with_imm_to_reg ),
//     .opcode_DIV_acc_by_reg_mem ( opcode_DIV_acc_by_reg_mem ),
//     .opcode_IDIV_acc_by_reg_mem ( opcode_IDIV_acc_by_reg_mem ),
//     .opcode_AAD ( opcode_AAD ),
//     .opcode_AAM ( opcode_AAM ),
//     .opcode_CBW ( opcode_CBW ),
//     .opcode_CWD ( opcode_CWD ),
//     .opcode_ROL_reg_mem_by_1 ( opcode_ROL_reg_mem_by_1 ),
//     .opcode_ROL_reg_mem_by_CL ( opcode_ROL_reg_mem_by_CL ),
//     .opcode_ROL_reg_mem_by_imm ( opcode_ROL_reg_mem_by_imm ),
//     .opcode_ROR_reg_mem_by_1 ( opcode_ROR_reg_mem_by_1 ),
//     .opcode_ROR_reg_mem_by_CL ( opcode_ROR_reg_mem_by_CL ),
//     .opcode_ROR_reg_mem_by_imm ( opcode_ROR_reg_mem_by_imm ),
//     .opcode_SHL_reg_mem_by_1 ( opcode_SHL_reg_mem_by_1 ),
//     .opcode_SHL_reg_mem_by_CL ( opcode_SHL_reg_mem_by_CL ),
//     .opcode_SHL_reg_mem_by_imm ( opcode_SHL_reg_mem_by_imm ),
//     .opcode_SAR_reg_mem_by_1 ( opcode_SAR_reg_mem_by_1 ),
//     .opcode_SAR_reg_mem_by_CL ( opcode_SAR_reg_mem_by_CL ),
//     .opcode_SAR_reg_mem_by_imm ( opcode_SAR_reg_mem_by_imm ),
//     .opcode_SHR_reg_mem_by_1 ( opcode_SHR_reg_mem_by_1 ),
//     .opcode_SHR_reg_mem_by_CL ( opcode_SHR_reg_mem_by_CL ),
//     .opcode_SHR_reg_mem_by_imm ( opcode_SHR_reg_mem_by_imm ),
//     .opcode_RCL_reg_mem_by_1 ( opcode_RCL_reg_mem_by_1 ),
//     .opcode_RCL_reg_mem_by_CL ( opcode_RCL_reg_mem_by_CL ),
//     .opcode_RCL_reg_mem_by_imm ( opcode_RCL_reg_mem_by_imm ),
//     .opcode_RCR_reg_mem_by_1 ( opcode_RCR_reg_mem_by_1 ),
//     .opcode_RCR_reg_mem_by_CL ( opcode_RCR_reg_mem_by_CL ),
//     .opcode_RCR_reg_mem_by_imm ( opcode_RCR_reg_mem_by_imm ),
//     .opcode_SHLD_reg_mem_by_imm ( opcode_SHLD_reg_mem_by_imm ),
//     .opcode_SHLD_reg_mem_by_CL ( opcode_SHLD_reg_mem_by_CL ),
//     .opcode_SHRD_reg_mem_by_imm ( opcode_SHRD_reg_mem_by_imm ),
//     .opcode_SHRD_reg_mem_by_CL ( opcode_SHRD_reg_mem_by_CL ),
//     .opcode_AND_reg_to_mem ( opcode_AND_reg_to_mem ),
//     .opcode_AND_mem_to_reg ( opcode_AND_mem_to_reg ),
//     .opcode_AND_imm_to_reg_mem ( opcode_AND_imm_to_reg_mem ),
//     .opcode_AND_imm_to_acc ( opcode_AND_imm_to_acc ),
//     .opcode_TEST_reg_mem_and_reg ( opcode_TEST_reg_mem_and_reg ),
//     .opcode_TEST_imm_to_reg_mem ( opcode_TEST_imm_to_reg_mem ),
//     .opcode_TEST_imm_to_acc ( opcode_TEST_imm_to_acc ),
//     .opcode_OR_reg_to_mem ( opcode_OR_reg_to_mem ),
//     .opcode_OR_mem_to_reg ( opcode_OR_mem_to_reg ),
//     .opcode_OR_imm_to_reg_mem ( opcode_OR_imm_to_reg_mem ),
//     .opcode_OR_imm_to_acc ( opcode_OR_imm_to_acc ),
//     .opcode_XOR_reg_to_mem ( opcode_XOR_reg_to_mem ),
//     .opcode_XOR_mem_to_reg ( opcode_XOR_mem_to_reg ),
//     .opcode_XOR_imm_to_reg_mem ( opcode_XOR_imm_to_reg_mem ),
//     .opcode_XOR_imm_to_acc ( opcode_XOR_imm_to_acc ),
//     .opcode_NOT ( opcode_NOT ),
//     .opcode_CMPS ( opcode_CMPS ),
//     .opcode_INS ( opcode_INS ),
//     .opcode_LODS ( opcode_LODS ),
//     .opcode_MOVS ( opcode_MOVS ),
//     .opcode_OUTS ( opcode_OUTS ),
//     .opcode_SCAS ( opcode_SCAS ),
//     .opcode_STOS ( opcode_STOS ),
//     .opcode_XLAT ( opcode_XLAT ),
//     .opcode_REPE ( opcode_REPE ),
//     .opcode_REPNE ( opcode_REPNE ),
//     .opcode_BSF ( opcode_BSF ),
//     .opcode_BSR ( opcode_BSR ),
//     .opcode_BT_reg_mem_with_imm ( opcode_BT_reg_mem_with_imm ),
//     .opcode_BT_reg_mem_with_reg ( opcode_BT_reg_mem_with_reg ),
//     .opcode_BTC_reg_mem_with_imm ( opcode_BTC_reg_mem_with_imm ),
//     .opcode_BTC_reg_mem_with_reg ( opcode_BTC_reg_mem_with_reg ),
//     .opcode_BTR_reg_mem_with_imm ( opcode_BTR_reg_mem_with_imm ),
//     .opcode_BTR_reg_mem_with_reg ( opcode_BTR_reg_mem_with_reg ),
//     .opcode_BTS_reg_mem_with_imm ( opcode_BTS_reg_mem_with_imm ),
//     .opcode_BTS_reg_mem_with_reg ( opcode_BTS_reg_mem_with_reg ),
//     .opcode_CALL_direct_within_segment ( opcode_CALL_direct_within_segment ),
//     .opcode_CALL_indirect_within_segment ( opcode_CALL_indirect_within_segment ),
//     .opcode_CALL_direct_intersegment ( opcode_CALL_direct_intersegment ),
//     .opcode_CALL_indirect_intersegment ( opcode_CALL_indirect_intersegment ),
//     .opcode_JMP_short ( opcode_JMP_short ),
//     .opcode_JMP_direct_within_segment ( opcode_JMP_direct_within_segment ),
//     .opcode_JMP_indirect_within_segment ( opcode_JMP_indirect_within_segment ),
//     .opcode_JMP_direct_intersegment ( opcode_JMP_direct_intersegment ),
//     .opcode_JMP_indirect_intersegment ( opcode_JMP_indirect_intersegment ),
//     .opcode_RET_within_segment ( opcode_RET_within_segment ),
//     .opcode_RET_within_segment_adding_imm_to_SP ( opcode_RET_within_segment_adding_imm_to_SP ),
//     .opcode_RET_intersegment ( opcode_RET_intersegment ),
//     .opcode_RET_intersegment_adding_imm_to_SP ( opcode_RET_intersegment_adding_imm_to_SP ),
//     .opcode_JO_8bit_disp ( opcode_JO_8bit_disp ),
//     .opcode_JO_full_disp ( opcode_JO_full_disp ),
//     .opcode_JNO_8bit_disp ( opcode_JNO_8bit_disp ),
//     .opcode_JNO_full_disp ( opcode_JNO_full_disp ),
//     .opcode_JB_8bit_disp ( opcode_JB_8bit_disp ),
//     .opcode_JB_full_disp ( opcode_JB_full_disp ),
//     .opcode_JNB_8bit_disp ( opcode_JNB_8bit_disp ),
//     .opcode_JNB_full_disp ( opcode_JNB_full_disp ),
//     .opcode_JE_8bit_disp ( opcode_JE_8bit_disp ),
//     .opcode_JE_full_disp ( opcode_JE_full_disp ),
//     .opcode_JNE_8bit_disp ( opcode_JNE_8bit_disp ),
//     .opcode_JNE_full_disp ( opcode_JNE_full_disp ),
//     .opcode_JBE_8bit_disp ( opcode_JBE_8bit_disp ),
//     .opcode_JBE_full_disp ( opcode_JBE_full_disp ),
//     .opcode_JNBE_8bit_disp ( opcode_JNBE_8bit_disp ),
//     .opcode_JNBE_full_disp ( opcode_JNBE_full_disp ),
//     .opcode_JS_8bit_disp ( opcode_JS_8bit_disp ),
//     .opcode_JS_full_disp ( opcode_JS_full_disp ),
//     .opcode_JNS_8bit_disp ( opcode_JNS_8bit_disp ),
//     .opcode_JNS_full_disp ( opcode_JNS_full_disp ),
//     .opcode_JP_8bit_disp ( opcode_JP_8bit_disp ),
//     .opcode_JP_full_disp ( opcode_JP_full_disp ),
//     .opcode_JNP_8bit_disp ( opcode_JNP_8bit_disp ),
//     .opcode_JNP_full_disp ( opcode_JNP_full_disp ),
//     .opcode_JL_8bit_disp ( opcode_JL_8bit_disp ),
//     .opcode_JL_full_disp ( opcode_JL_full_disp ),
//     .opcode_JNL_8bit_disp ( opcode_JNL_8bit_disp ),
//     .opcode_JNL_full_disp ( opcode_JNL_full_disp ),
//     .opcode_JLE_8bit_disp ( opcode_JLE_8bit_disp ),
//     .opcode_JLE_full_disp ( opcode_JLE_full_disp ),
//     .opcode_JNLE_8bit_disp ( opcode_JNLE_8bit_disp ),
//     .opcode_JNLE_full_disp ( opcode_JNLE_full_disp ),
//     .opcode_JCXZ ( opcode_JCXZ ),
//     .opcode_LOOP ( opcode_LOOP ),
//     .opcode_LOOPZ ( opcode_LOOPZ ),
//     .opcode_LOOPNZ ( opcode_LOOPNZ ),
//     .opcode_SETO ( opcode_SETO ),
//     .opcode_SETNO ( opcode_SETNO ),
//     .opcode_SETB ( opcode_SETB ),
//     .opcode_SETNB ( opcode_SETNB ),
//     .opcode_SETE ( opcode_SETE ),
//     .opcode_SETNE ( opcode_SETNE ),
//     .opcode_SETBE ( opcode_SETBE ),
//     .opcode_SETNBE ( opcode_SETNBE ),
//     .opcode_SETS ( opcode_SETS ),
//     .opcode_SETNS ( opcode_SETNS ),
//     .opcode_SETP ( opcode_SETP ),
//     .opcode_SETNP ( opcode_SETNP ),
//     .opcode_SETL ( opcode_SETL ),
//     .opcode_SETNL ( opcode_SETNL ),
//     .opcode_SETLE ( opcode_SETLE ),
//     .opcode_SETNLE ( opcode_SETNLE ),
//     .opcode_ENTER ( opcode_ENTER ),
//     .opcode_LEAVE ( opcode_LEAVE ),
//     .opcode_INT_type_3 ( opcode_INT_type_3 ),
//     .opcode_INT_type_specified ( opcode_INT_type_specified ),
//     .opcode_INTO ( opcode_INTO ),
//     .opcode_BOUND ( opcode_BOUND ),
//     .opcode_IRET ( opcode_IRET ),
//     .opcode_HLT ( opcode_HLT ),
//     .opcode_MOV_CR0_CR2_CR3_from_reg ( opcode_MOV_CR0_CR2_CR3_from_reg ),
//     .opcode_MOV_reg_from_CR0_3 ( opcode_MOV_reg_from_CR0_3 ),
//     .opcode_MOV_DR0_7_from_reg ( opcode_MOV_DR0_7_from_reg ),
//     .opcode_MOV_reg_from_DR0_7 ( opcode_MOV_reg_from_DR0_7 ),
//     .opcode_MOV_TR6_7_from_reg ( opcode_MOV_TR6_7_from_reg ),
//     .opcode_MOV_reg_from_TR6_7 ( opcode_MOV_reg_from_TR6_7 ),
//     .opcode_NOP ( opcode_NOP ),
//     .opcode_WAIT ( opcode_WAIT ),
//     .opcode_processor_extension_escape ( opcode_processor_extension_escape ),
//     .opcode_prefix_address_size ( opcode_prefix_address_size ),
//     .opcode_prefix_bus_lock ( opcode_prefix_bus_lock ),
//     .opcode_prefix_operand_size ( opcode_prefix_operand_size ),
//     .opcode_prefix_segment_override_CS ( opcode_prefix_segment_override_CS ),
//     .opcode_prefix_segment_override_DS ( opcode_prefix_segment_override_DS ),
//     .opcode_prefix_segment_override_ES ( opcode_prefix_segment_override_ES ),
//     .opcode_prefix_segment_override_FS ( opcode_prefix_segment_override_FS ),
//     .opcode_prefix_segment_override_GS ( opcode_prefix_segment_override_GS ),
//     .opcode_prefix_segment_override_SS ( opcode_prefix_segment_override_SS ),
//     .opcode_ARPL ( opcode_ARPL ),
//     .opcode_LAR ( opcode_LAR ),
//     .opcode_LGDT ( opcode_LGDT ),
//     .opcode_LIDT ( opcode_LIDT ),
//     .opcode_LLDT ( opcode_LLDT ),
//     .opcode_LMSW ( opcode_LMSW ),
//     .opcode_LSL ( opcode_LSL ),
//     .opcode_LTR ( opcode_LTR ),
//     .opcode_SGDT ( opcode_SGDT ),
//     .opcode_SIDT ( opcode_SIDT ),
//     .opcode_SLDT ( opcode_SLDT ),
//     .opcode_SMSW ( opcode_SMSW ),
//     .opcode_STR ( opcode_STR ),
//     .opcode_VERR ( opcode_VERR ),
//     .opcode_VERW ( opcode_VERW ),
//     .instruction ( instruction ),
//     .s ( s ),
//     .w ( w ),
//     .gereral_propose_register ( gereral_propose_register ),
//     .sreg ( sreg ),
//     .mod ( mod ),
//     .rm ( rm ),
//     .has_s ( has_s ),
//     .has_w ( has_w ),
//     .has_sreg ( has_sreg ),
//     .has_mod_rm ( has_mod_rm ),
//     .is_prefix_segment ( is_prefix_segment ),
//     .is_prefix ( is_prefix )
// );

// logic length_1;
// logic length_2;
// logic length_3;
// logic length_4;
// decode_opcode_length u_decode_opcode_length (
//     .opcode_MOV_reg_to_reg_mem ( opcode_MOV_reg_to_reg_mem ),
//     .opcode_MOV_reg_mem_to_reg ( opcode_MOV_reg_mem_to_reg ),
//     .opcode_MOV_imm_to_reg_mem ( opcode_MOV_imm_to_reg_mem ),
//     .opcode_MOV_imm_to_reg_short ( opcode_MOV_imm_to_reg_short ),
//     .opcode_MOV_mem_to_acc ( opcode_MOV_mem_to_acc ),
//     .opcode_MOV_acc_to_mem ( opcode_MOV_acc_to_mem ),
//     .opcode_MOV_reg_mem_to_sreg ( opcode_MOV_reg_mem_to_sreg ),
//     .opcode_MOV_sreg_to_reg_mem ( opcode_MOV_sreg_to_reg_mem ),
//     .opcode_MOVSX ( opcode_MOVSX ),
//     .opcode_MOVZX ( opcode_MOVZX ),
//     .opcode_PUSH_reg_mem ( opcode_PUSH_reg_mem ),
//     .opcode_PUSH_reg_short ( opcode_PUSH_reg_short ),
//     .opcode_PUSH_sreg_2 ( opcode_PUSH_sreg_2 ),
//     .opcode_PUSH_sreg_3 ( opcode_PUSH_sreg_3 ),
//     .opcode_PUSH_imm ( opcode_PUSH_imm ),
//     .opcode_PUSH_all ( opcode_PUSH_all ),
//     .opcode_POP_reg_mem ( opcode_POP_reg_mem ),
//     .opcode_POP_reg_short ( opcode_POP_reg_short ),
//     .opcode_POP_sreg_2 ( opcode_POP_sreg_2 ),
//     .opcode_POP_sreg_3 ( opcode_POP_sreg_3 ),
//     .opcode_POP_all ( opcode_POP_all ),
//     .opcode_XCHG_reg_mem_with_reg ( opcode_XCHG_reg_mem_with_reg ),
//     .opcode_XCHG_reg_with_acc_short ( opcode_XCHG_reg_with_acc_short ),
//     .opcode_IN_port_fixed ( opcode_IN_port_fixed ),
//     .opcode_IN_port_variable ( opcode_IN_port_variable ),
//     .opcode_OUT_port_fixed ( opcode_OUT_port_fixed ),
//     .opcode_OUT_port_variable ( opcode_OUT_port_variable ),
//     .opcode_LEA_load_ea_to_reg ( opcode_LEA_load_ea_to_reg ),
//     .opcode_LDS_load_ptr_to_DS ( opcode_LDS_load_ptr_to_DS ),
//     .opcode_LES_load_ptr_to_ES ( opcode_LES_load_ptr_to_ES ),
//     .opcode_LFS_load_ptr_to_FS ( opcode_LFS_load_ptr_to_FS ),
//     .opcode_LGS_load_ptr_to_GS ( opcode_LGS_load_ptr_to_GS ),
//     .opcode_LSS_load_ptr_to_SS ( opcode_LSS_load_ptr_to_SS ),
//     .opcode_CLC_clear_carry_flag ( opcode_CLC_clear_carry_flag ),
//     .opcode_CLD_clear_direction_flag ( opcode_CLD_clear_direction_flag ),
//     .opcode_CLI_clear_interrupt_enable_flag ( opcode_CLI_clear_interrupt_enable_flag ),
//     .opcode_CLTS_clear_task_switched_flag ( opcode_CLTS_clear_task_switched_flag ),
//     .opcode_CMC_complement_carry_flag ( opcode_CMC_complement_carry_flag ),
//     .opcode_LAHF_load_ah_into_flag ( opcode_LAHF_load_ah_into_flag ),
//     .opcode_POPF_pop_flags ( opcode_POPF_pop_flags ),
//     .opcode_PUSHF_push_flags ( opcode_PUSHF_push_flags ),
//     .opcode_SAHF_store_ah_into_flag ( opcode_SAHF_store_ah_into_flag ),
//     .opcode_STC_set_carry_flag ( opcode_STC_set_carry_flag ),
//     .opcode_STD_set_direction_flag ( opcode_STD_set_direction_flag ),
//     .opcode_STI_set_interrupt_enable_flag ( opcode_STI_set_interrupt_enable_flag ),
//     .opcode_ADD_reg_to_mem ( opcode_ADD_reg_to_mem ),
//     .opcode_ADD_mem_to_reg ( opcode_ADD_mem_to_reg ),
//     .opcode_ADD_imm_to_reg_mem ( opcode_ADD_imm_to_reg_mem ),
//     .opcode_ADD_imm_to_acc ( opcode_ADD_imm_to_acc ),
//     .opcode_ADC_reg_to_mem ( opcode_ADC_reg_to_mem ),
//     .opcode_ADC_mem_to_reg ( opcode_ADC_mem_to_reg ),
//     .opcode_ADC_imm_to_reg_mem ( opcode_ADC_imm_to_reg_mem ),
//     .opcode_ADC_imm_to_acc ( opcode_ADC_imm_to_acc ),
//     .opcode_INC_reg_mem ( opcode_INC_reg_mem ),
//     .opcode_INC_reg ( opcode_INC_reg ),
//     .opcode_SUB_reg_to_mem ( opcode_SUB_reg_to_mem ),
//     .opcode_SUB_mem_to_reg ( opcode_SUB_mem_to_reg ),
//     .opcode_SUB_imm_to_reg_mem ( opcode_SUB_imm_to_reg_mem ),
//     .opcode_SUB_imm_to_acc ( opcode_SUB_imm_to_acc ),
//     .opcode_SBB_reg_to_mem ( opcode_SBB_reg_to_mem ),
//     .opcode_SBB_mem_to_reg ( opcode_SBB_mem_to_reg ),
//     .opcode_SBB_imm_to_reg_mem ( opcode_SBB_imm_to_reg_mem ),
//     .opcode_SBB_imm_to_acc ( opcode_SBB_imm_to_acc ),
//     .opcode_DEC_reg_mem ( opcode_DEC_reg_mem ),
//     .opcode_DEC_reg ( opcode_DEC_reg ),
//     .opcode_CMP_mem_with_reg ( opcode_CMP_mem_with_reg ),
//     .opcode_CMP_reg_with_mem ( opcode_CMP_reg_with_mem ),
//     .opcode_CMP_imm_with_reg_mem ( opcode_CMP_imm_with_reg_mem ),
//     .opcode_CMP_imm_with_acc ( opcode_CMP_imm_with_acc ),
//     .opcode_NEG_change_sign ( opcode_NEG_change_sign ),
//     .opcode_AAA ( opcode_AAA ),
//     .opcode_AAS ( opcode_AAS ),
//     .opcode_DAA ( opcode_DAA ),
//     .opcode_DAS ( opcode_DAS ),
//     .opcode_MUL_acc_with_reg_mem ( opcode_MUL_acc_with_reg_mem ),
//     .opcode_IMUL_acc_with_reg_mem ( opcode_IMUL_acc_with_reg_mem ),
//     .opcode_IMUL_reg_with_reg_mem ( opcode_IMUL_reg_with_reg_mem ),
//     .opcode_IMUL_reg_mem_with_imm_to_reg ( opcode_IMUL_reg_mem_with_imm_to_reg ),
//     .opcode_DIV_acc_by_reg_mem ( opcode_DIV_acc_by_reg_mem ),
//     .opcode_IDIV_acc_by_reg_mem ( opcode_IDIV_acc_by_reg_mem ),
//     .opcode_AAD ( opcode_AAD ),
//     .opcode_AAM ( opcode_AAM ),
//     .opcode_CBW ( opcode_CBW ),
//     .opcode_CWD ( opcode_CWD ),
//     .opcode_ROL_reg_mem_by_1 ( opcode_ROL_reg_mem_by_1 ),
//     .opcode_ROL_reg_mem_by_CL ( opcode_ROL_reg_mem_by_CL ),
//     .opcode_ROL_reg_mem_by_imm ( opcode_ROL_reg_mem_by_imm ),
//     .opcode_ROR_reg_mem_by_1 ( opcode_ROR_reg_mem_by_1 ),
//     .opcode_ROR_reg_mem_by_CL ( opcode_ROR_reg_mem_by_CL ),
//     .opcode_ROR_reg_mem_by_imm ( opcode_ROR_reg_mem_by_imm ),
//     .opcode_SHL_reg_mem_by_1 ( opcode_SHL_reg_mem_by_1 ),
//     .opcode_SHL_reg_mem_by_CL ( opcode_SHL_reg_mem_by_CL ),
//     .opcode_SHL_reg_mem_by_imm ( opcode_SHL_reg_mem_by_imm ),
//     .opcode_SAR_reg_mem_by_1 ( opcode_SAR_reg_mem_by_1 ),
//     .opcode_SAR_reg_mem_by_CL ( opcode_SAR_reg_mem_by_CL ),
//     .opcode_SAR_reg_mem_by_imm ( opcode_SAR_reg_mem_by_imm ),
//     .opcode_SHR_reg_mem_by_1 ( opcode_SHR_reg_mem_by_1 ),
//     .opcode_SHR_reg_mem_by_CL ( opcode_SHR_reg_mem_by_CL ),
//     .opcode_SHR_reg_mem_by_imm ( opcode_SHR_reg_mem_by_imm ),
//     .opcode_RCL_reg_mem_by_1 ( opcode_RCL_reg_mem_by_1 ),
//     .opcode_RCL_reg_mem_by_CL ( opcode_RCL_reg_mem_by_CL ),
//     .opcode_RCL_reg_mem_by_imm ( opcode_RCL_reg_mem_by_imm ),
//     .opcode_RCR_reg_mem_by_1 ( opcode_RCR_reg_mem_by_1 ),
//     .opcode_RCR_reg_mem_by_CL ( opcode_RCR_reg_mem_by_CL ),
//     .opcode_RCR_reg_mem_by_imm ( opcode_RCR_reg_mem_by_imm ),
//     .opcode_SHLD_reg_mem_by_imm ( opcode_SHLD_reg_mem_by_imm ),
//     .opcode_SHLD_reg_mem_by_CL ( opcode_SHLD_reg_mem_by_CL ),
//     .opcode_SHRD_reg_mem_by_imm ( opcode_SHRD_reg_mem_by_imm ),
//     .opcode_SHRD_reg_mem_by_CL ( opcode_SHRD_reg_mem_by_CL ),
//     .opcode_AND_reg_to_mem ( opcode_AND_reg_to_mem ),
//     .opcode_AND_mem_to_reg ( opcode_AND_mem_to_reg ),
//     .opcode_AND_imm_to_reg_mem ( opcode_AND_imm_to_reg_mem ),
//     .opcode_AND_imm_to_acc ( opcode_AND_imm_to_acc ),
//     .opcode_TEST_reg_mem_and_reg ( opcode_TEST_reg_mem_and_reg ),
//     .opcode_TEST_imm_to_reg_mem ( opcode_TEST_imm_to_reg_mem ),
//     .opcode_TEST_imm_to_acc ( opcode_TEST_imm_to_acc ),
//     .opcode_OR_reg_to_mem ( opcode_OR_reg_to_mem ),
//     .opcode_OR_mem_to_reg ( opcode_OR_mem_to_reg ),
//     .opcode_OR_imm_to_reg_mem ( opcode_OR_imm_to_reg_mem ),
//     .opcode_OR_imm_to_acc ( opcode_OR_imm_to_acc ),
//     .opcode_XOR_reg_to_mem ( opcode_XOR_reg_to_mem ),
//     .opcode_XOR_mem_to_reg ( opcode_XOR_mem_to_reg ),
//     .opcode_XOR_imm_to_reg_mem ( opcode_XOR_imm_to_reg_mem ),
//     .opcode_XOR_imm_to_acc ( opcode_XOR_imm_to_acc ),
//     .opcode_NOT ( opcode_NOT ),
//     .opcode_CMPS ( opcode_CMPS ),
//     .opcode_INS ( opcode_INS ),
//     .opcode_LODS ( opcode_LODS ),
//     .opcode_MOVS ( opcode_MOVS ),
//     .opcode_OUTS ( opcode_OUTS ),
//     .opcode_SCAS ( opcode_SCAS ),
//     .opcode_STOS ( opcode_STOS ),
//     .opcode_XLAT ( opcode_XLAT ),
//     .opcode_REPE ( opcode_REPE ),
//     .opcode_REPNE ( opcode_REPNE ),
//     .opcode_BSF ( opcode_BSF ),
//     .opcode_BSR ( opcode_BSR ),
//     .opcode_BT_reg_mem_with_imm ( opcode_BT_reg_mem_with_imm ),
//     .opcode_BT_reg_mem_with_reg ( opcode_BT_reg_mem_with_reg ),
//     .opcode_BTC_reg_mem_with_imm ( opcode_BTC_reg_mem_with_imm ),
//     .opcode_BTC_reg_mem_with_reg ( opcode_BTC_reg_mem_with_reg ),
//     .opcode_BTR_reg_mem_with_imm ( opcode_BTR_reg_mem_with_imm ),
//     .opcode_BTR_reg_mem_with_reg ( opcode_BTR_reg_mem_with_reg ),
//     .opcode_BTS_reg_mem_with_imm ( opcode_BTS_reg_mem_with_imm ),
//     .opcode_BTS_reg_mem_with_reg ( opcode_BTS_reg_mem_with_reg ),
//     .opcode_CALL_direct_within_segment ( opcode_CALL_direct_within_segment ),
//     .opcode_CALL_indirect_within_segment ( opcode_CALL_indirect_within_segment ),
//     .opcode_CALL_direct_intersegment ( opcode_CALL_direct_intersegment ),
//     .opcode_CALL_indirect_intersegment ( opcode_CALL_indirect_intersegment ),
//     .opcode_JMP_short ( opcode_JMP_short ),
//     .opcode_JMP_direct_within_segment ( opcode_JMP_direct_within_segment ),
//     .opcode_JMP_indirect_within_segment ( opcode_JMP_indirect_within_segment ),
//     .opcode_JMP_direct_intersegment ( opcode_JMP_direct_intersegment ),
//     .opcode_JMP_indirect_intersegment ( opcode_JMP_indirect_intersegment ),
//     .opcode_RET_within_segment ( opcode_RET_within_segment ),
//     .opcode_RET_within_segment_adding_imm_to_SP ( opcode_RET_within_segment_adding_imm_to_SP ),
//     .opcode_RET_intersegment ( opcode_RET_intersegment ),
//     .opcode_RET_intersegment_adding_imm_to_SP ( opcode_RET_intersegment_adding_imm_to_SP ),
//     .opcode_JO_8bit_disp ( opcode_JO_8bit_disp ),
//     .opcode_JO_full_disp ( opcode_JO_full_disp ),
//     .opcode_JNO_8bit_disp ( opcode_JNO_8bit_disp ),
//     .opcode_JNO_full_disp ( opcode_JNO_full_disp ),
//     .opcode_JB_8bit_disp ( opcode_JB_8bit_disp ),
//     .opcode_JB_full_disp ( opcode_JB_full_disp ),
//     .opcode_JNB_8bit_disp ( opcode_JNB_8bit_disp ),
//     .opcode_JNB_full_disp ( opcode_JNB_full_disp ),
//     .opcode_JE_8bit_disp ( opcode_JE_8bit_disp ),
//     .opcode_JE_full_disp ( opcode_JE_full_disp ),
//     .opcode_JNE_8bit_disp ( opcode_JNE_8bit_disp ),
//     .opcode_JNE_full_disp ( opcode_JNE_full_disp ),
//     .opcode_JBE_8bit_disp ( opcode_JBE_8bit_disp ),
//     .opcode_JBE_full_disp ( opcode_JBE_full_disp ),
//     .opcode_JNBE_8bit_disp ( opcode_JNBE_8bit_disp ),
//     .opcode_JNBE_full_disp ( opcode_JNBE_full_disp ),
//     .opcode_JS_8bit_disp ( opcode_JS_8bit_disp ),
//     .opcode_JS_full_disp ( opcode_JS_full_disp ),
//     .opcode_JNS_8bit_disp ( opcode_JNS_8bit_disp ),
//     .opcode_JNS_full_disp ( opcode_JNS_full_disp ),
//     .opcode_JP_8bit_disp ( opcode_JP_8bit_disp ),
//     .opcode_JP_full_disp ( opcode_JP_full_disp ),
//     .opcode_JNP_8bit_disp ( opcode_JNP_8bit_disp ),
//     .opcode_JNP_full_disp ( opcode_JNP_full_disp ),
//     .opcode_JL_8bit_disp ( opcode_JL_8bit_disp ),
//     .opcode_JL_full_disp ( opcode_JL_full_disp ),
//     .opcode_JNL_8bit_disp ( opcode_JNL_8bit_disp ),
//     .opcode_JNL_full_disp ( opcode_JNL_full_disp ),
//     .opcode_JLE_8bit_disp ( opcode_JLE_8bit_disp ),
//     .opcode_JLE_full_disp ( opcode_JLE_full_disp ),
//     .opcode_JNLE_8bit_disp ( opcode_JNLE_8bit_disp ),
//     .opcode_JNLE_full_disp ( opcode_JNLE_full_disp ),
//     .opcode_JCXZ ( opcode_JCXZ ),
//     .opcode_LOOP ( opcode_LOOP ),
//     .opcode_LOOPZ ( opcode_LOOPZ ),
//     .opcode_LOOPNZ ( opcode_LOOPNZ ),
//     .opcode_SETO ( opcode_SETO ),
//     .opcode_SETNO ( opcode_SETNO ),
//     .opcode_SETB ( opcode_SETB ),
//     .opcode_SETNB ( opcode_SETNB ),
//     .opcode_SETE ( opcode_SETE ),
//     .opcode_SETNE ( opcode_SETNE ),
//     .opcode_SETBE ( opcode_SETBE ),
//     .opcode_SETNBE ( opcode_SETNBE ),
//     .opcode_SETS ( opcode_SETS ),
//     .opcode_SETNS ( opcode_SETNS ),
//     .opcode_SETP ( opcode_SETP ),
//     .opcode_SETNP ( opcode_SETNP ),
//     .opcode_SETL ( opcode_SETL ),
//     .opcode_SETNL ( opcode_SETNL ),
//     .opcode_SETLE ( opcode_SETLE ),
//     .opcode_SETNLE ( opcode_SETNLE ),
//     .opcode_ENTER ( opcode_ENTER ),
//     .opcode_LEAVE ( opcode_LEAVE ),
//     .opcode_INT_type_3 ( opcode_INT_type_3 ),
//     .opcode_INT_type_specified ( opcode_INT_type_specified ),
//     .opcode_INTO ( opcode_INTO ),
//     .opcode_BOUND ( opcode_BOUND ),
//     .opcode_IRET ( opcode_IRET ),
//     .opcode_HLT ( opcode_HLT ),
//     .opcode_MOV_CR0_CR2_CR3_from_reg ( opcode_MOV_CR0_CR2_CR3_from_reg ),
//     .opcode_MOV_reg_from_CR0_3 ( opcode_MOV_reg_from_CR0_3 ),
//     .opcode_MOV_DR0_7_from_reg ( opcode_MOV_DR0_7_from_reg ),
//     .opcode_MOV_reg_from_DR0_7 ( opcode_MOV_reg_from_DR0_7 ),
//     .opcode_MOV_TR6_7_from_reg ( opcode_MOV_TR6_7_from_reg ),
//     .opcode_MOV_reg_from_TR6_7 ( opcode_MOV_reg_from_TR6_7 ),
//     .opcode_NOP ( opcode_NOP ),
//     .opcode_WAIT ( opcode_WAIT ),
//     .opcode_processor_extension_escape ( opcode_processor_extension_escape ),
//     .opcode_prefix_address_size ( opcode_prefix_address_size ),
//     .opcode_prefix_bus_lock ( opcode_prefix_bus_lock ),
//     .opcode_prefix_operand_size ( opcode_prefix_operand_size ),
//     .opcode_prefix_segment_override_CS ( opcode_prefix_segment_override_CS ),
//     .opcode_prefix_segment_override_DS ( opcode_prefix_segment_override_DS ),
//     .opcode_prefix_segment_override_ES ( opcode_prefix_segment_override_ES ),
//     .opcode_prefix_segment_override_FS ( opcode_prefix_segment_override_FS ),
//     .opcode_prefix_segment_override_GS ( opcode_prefix_segment_override_GS ),
//     .opcode_prefix_segment_override_SS ( opcode_prefix_segment_override_SS ),
//     .opcode_ARPL ( opcode_ARPL ),
//     .opcode_LAR ( opcode_LAR ),
//     .opcode_LGDT ( opcode_LGDT ),
//     .opcode_LIDT ( opcode_LIDT ),
//     .opcode_LLDT ( opcode_LLDT ),
//     .opcode_LMSW ( opcode_LMSW ),
//     .opcode_LSL ( opcode_LSL ),
//     .opcode_LTR ( opcode_LTR ),
//     .opcode_SGDT ( opcode_SGDT ),
//     .opcode_SIDT ( opcode_SIDT ),
//     .opcode_SLDT ( opcode_SLDT ),
//     .opcode_SMSW ( opcode_SMSW ),
//     .opcode_STR ( opcode_STR ),
//     .opcode_VERR ( opcode_VERR ),
//     .opcode_VERW ( opcode_VERW ),
//     .length_1 ( length_1 ),
//     .length_2 ( length_2 ),
//     .length_3 ( length_3 ),
//     .length_4 ( length_4 )
// );

// decode_mod_rm u_decode_mod_rm (
//     .mod ( mod ),
//     .rm ( rm ),
//     .w ( w ),
//     .info_bit_width ( bit_width ),
//     .info_segment_reg ( info_segment_reg ),
//     .info_base_reg ( info_base_reg ),
//     .info_index_reg ( info_index_reg ),
//     .info_displacement ( info_displacement ),
//     .sib_is_present ( sib_is_present )
// );


endmodule
