module soc_top (
    input  logic        clock,
    input  logic        reset
);

w80386_cpu cpu_0 ();

/*
connect to:
RAM
BIOS ROM
VGA
PS/2 mouse and keyboard
Audio
Ethernet
*/

endmodule