/*
project: w80386dx
author: Chang Wei<changwei1006@gmail.com>
repo: https://github.com/openx86/w80386dx
module: decode unit
create at: 2022-01-04 03:27:51
description: decode unit module
*/

`include "D:/GitHub/openx86/w80386dx/rtl/definition.h"

module decode (
    input  logic [ 7:0] i_instruction [0:15],
    input  logic        i_default_operand_size,
    output logic        o_group_1_lock_bus,
    output logic        o_group_1_repeat_not_equal,
    output logic        o_group_1_repeat_equal,
    output logic        o_group_1_bound,
    output logic        o_group_2_segment_override,
    output logic        o_group_2_hint_branch_not_taken,
    output logic        o_group_2_hint_branch_taken,
    output logic        o_group_3_operand_size,
    output logic        o_group_4_address_size,
    output logic [ 2:0] o_segment_override_index,
    output logic        o_consume_bytes_prefix_1,
    output logic        o_consume_bytes_prefix_2,
    output logic        o_consume_bytes_prefix_3,
    output logic        o_consume_bytes_prefix_4,
    output logic        o_error_stage_1,
    output logic        o_x86_ADC_reg_1_to_reg_2,
    output logic        o_x86_ADC_reg_2_to_reg_1,
    output logic        o_x86_ADC_mem_to_reg,
    output logic        o_x86_ADC_reg_to_mem,
    output logic        o_x86_ADC_imm_to_reg,
    output logic        o_x86_ADC_imm_to_acc,
    output logic        o_x86_ADC_imm_to_mem,
    output logic        o_error_stage_2,
    output logic [ 2:0] o_index_reg_gen [0:2],
    output logic        o_index_reg_gen_is_present,
    output logic [ 2:0] o_index_reg_seg,
    output logic        o_index_reg_seg_is_present,
    output logic        o_w_is_present,
    output logic        o_w,
    output logic        o_s_is_present,
    output logic        o_s,
    output logic        o_mod_rm_is_present,
    output logic [ 1:0] o_mod,
    output logic [ 2:0] o_rm,
    output logic        o_immediate_size_f,
    output logic        o_consume_bytes_opcode_1,
    output logic        o_consume_bytes_opcode_2,
    output logic        o_consume_bytes_opcode_3,
    output logic        o_error_stage_3,
    output logic [ 2:0] o_segment_reg_index,
    output logic        o_base_reg_is_present,
    output logic [ 2:0] o_base_reg_index,
    output logic        o_index_reg_is_present,
    output logic [ 2:0] o_index_reg_index,
    output logic        o_displacement_size_1,
    output logic        o_displacement_size_2,
    output logic        o_displacement_size_4,
    output logic        o_sib_is_present,
    output logic [ 1:0] o_scale_factor,
    output logic        o_error_stage_4,
    output logic [31:0] o_displacement,
    output logic [31:0] o_immediate,
    output logic [ 3:0] o_consume_bytes,
    output logic        o_error_stage_5,

    // output logic [ 2:0] o_index_reg_gen [0:2],
    // output logic [ 2:0] o_index_reg_seg,
    // output logic [ 2:0] o_index_reg_base,
    // output logic [ 2:0] o_index_reg_index,
    // output logic [ 1:0] o_index_scale_factor,
    // output logic [31:0] o_displacement,
    // output logic [31:0] o_immediate,
    output logic        o_error
);

decode_stage_1 (
    i_instruction,
    i_default_operand_size,
    o_group_1_lock_bus,
    o_group_1_repeat_not_equal,
    o_group_1_repeat_equal,
    o_group_1_bound,
    o_group_2_segment_override,
    o_group_2_hint_branch_not_taken,
    o_group_2_hint_branch_taken,
    o_group_3_operand_size,
    o_group_4_address_size,
    o_segment_override_index,
    o_consume_bytes_prefix_1,
    o_consume_bytes_prefix_2,
    o_consume_bytes_prefix_3,
    o_consume_bytes_prefix_4,
    o_error_stage_1
);

decode_stage_2 (
    i_instruction,
    i_default_operand_size,
    o_group_1_lock_bus,
    o_group_1_repeat_not_equal,
    o_group_1_repeat_equal,
    o_group_1_bound,
    o_group_2_segment_override,
    o_group_2_hint_branch_not_taken,
    o_group_2_hint_branch_taken,
    o_group_3_operand_size,
    o_group_4_address_size,
    o_segment_override_index,
    o_consume_bytes_prefix_1,
    o_consume_bytes_prefix_2,
    o_consume_bytes_prefix_3,
    o_consume_bytes_prefix_4,
    o_error_stage_1,
    o_x86_ADC_reg_1_to_reg_2,
    o_x86_ADC_reg_2_to_reg_1,
    o_x86_ADC_mem_to_reg,
    o_x86_ADC_reg_to_mem,
    o_x86_ADC_imm_to_reg,
    o_x86_ADC_imm_to_acc,
    o_x86_ADC_imm_to_mem,
    o_error_stage_2
);

decode_stage_3 (
    i_instruction,
    i_default_operand_size,
    o_group_1_lock_bus,
    o_group_1_repeat_not_equal,
    o_group_1_repeat_equal,
    o_group_1_bound,
    o_group_2_segment_override,
    o_group_2_hint_branch_not_taken,
    o_group_2_hint_branch_taken,
    o_group_3_operand_size,
    o_group_4_address_size,
    o_segment_override_index,
    o_consume_bytes_prefix_1,
    o_consume_bytes_prefix_2,
    o_consume_bytes_prefix_3,
    o_consume_bytes_prefix_4,
    o_error_stage_1,
    o_x86_ADC_reg_1_to_reg_2,
    o_x86_ADC_reg_2_to_reg_1,
    o_x86_ADC_mem_to_reg,
    o_x86_ADC_reg_to_mem,
    o_x86_ADC_imm_to_reg,
    o_x86_ADC_imm_to_acc,
    o_x86_ADC_imm_to_mem,
    o_error_stage_2,
    o_index_reg_gen,
    o_index_reg_gen_is_present,
    o_index_reg_seg,
    o_index_reg_seg_is_present,
    o_w_is_present,
    o_w,
    o_s_is_present,
    o_s,
    o_mod_rm_is_present,
    o_mod,
    o_rm,
    o_immediate_size_full,
    o_consume_bytes_opcode_1,
    o_consume_bytes_opcode_2,
    o_consume_bytes_opcode_3,
    o_error_stage_3
);

decode_stage_4 (
    i_instruction,
    i_default_operand_size,
    o_group_1_lock_bus,
    o_group_1_repeat_not_equal,
    o_group_1_repeat_equal,
    o_group_1_bound,
    o_group_2_segment_override,
    o_group_2_hint_branch_not_taken,
    o_group_2_hint_branch_taken,
    o_group_3_operand_size,
    o_group_4_address_size,
    o_segment_override_index,
    o_consume_bytes_prefix_1,
    o_consume_bytes_prefix_2,
    o_consume_bytes_prefix_3,
    o_consume_bytes_prefix_4,
    o_error_stage_1,
    o_x86_ADC_reg_1_to_reg_2,
    o_x86_ADC_reg_2_to_reg_1,
    o_x86_ADC_mem_to_reg,
    o_x86_ADC_reg_to_mem,
    o_x86_ADC_imm_to_reg,
    o_x86_ADC_imm_to_acc,
    o_x86_ADC_imm_to_mem,
    o_error_stage_2,
    o_index_reg_gen,
    o_index_reg_gen_is_present,
    o_index_reg_seg,
    o_index_reg_seg_is_present,
    o_w_is_present,
    o_w,
    o_s_is_present,
    o_s,
    o_mod_rm_is_present,
    o_mod,
    o_rm,
    o_immediate_size_full,
    o_consume_bytes_opcode_1,
    o_consume_bytes_opcode_2,
    o_consume_bytes_opcode_3,
    o_error_stage_3,
    o_segment_reg_index,
    o_base_reg_is_present,
    o_base_reg_index,
    o_index_reg_is_present,
    o_index_reg_index,
    o_displacement_size_1,
    o_displacement_size_2,
    o_displacement_size_4,
    o_scale_factor,
    o_error_stage_4
);

decode_stage_5 (
    i_instruction,
    i_default_operand_size,
    o_group_1_lock_bus,
    o_group_1_repeat_not_equal,
    o_group_1_repeat_equal,
    o_group_1_bound,
    o_group_2_segment_override,
    o_group_2_hint_branch_not_taken,
    o_group_2_hint_branch_taken,
    o_group_3_operand_size,
    o_group_4_address_size,
    o_segment_override_index,
    o_consume_bytes_prefix_1,
    o_consume_bytes_prefix_2,
    o_consume_bytes_prefix_3,
    o_consume_bytes_prefix_4,
    o_error_stage_1,
    o_x86_ADC_reg_1_to_reg_2,
    o_x86_ADC_reg_2_to_reg_1,
    o_x86_ADC_mem_to_reg,
    o_x86_ADC_reg_to_mem,
    o_x86_ADC_imm_to_reg,
    o_x86_ADC_imm_to_acc,
    o_x86_ADC_imm_to_mem,
    o_error_stage_2,
    o_index_reg_gen,
    o_index_reg_gen_is_present,
    o_index_reg_seg,
    o_index_reg_seg_is_present,
    o_w_is_present,
    o_w,
    o_s_is_present,
    o_s,
    o_mod_rm_is_present,
    o_mod,
    o_rm,
    o_immediate_size_full,
    o_consume_bytes_opcode_1,
    o_consume_bytes_opcode_2,
    o_consume_bytes_opcode_3,
    o_error_stage_3,
    o_segment_reg_index,
    o_base_reg_is_present,
    o_base_reg_index,
    o_index_reg_is_present,
    o_index_reg_index,
    o_displacement_size_1,
    o_displacement_size_2,
    o_displacement_size_4,
    o_scale_factor,
    o_error_stage_4,
    o_displacement,
    o_immediate,
    o_consume_bytes,
    o_error_stage_5
);

endmodule
