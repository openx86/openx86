/*
project: w80386dx
author: Chang Wei<changwei1006@gmail.com>
repo: https://github.com/openx86/w80386dx
module: decode_field
create at: 2021-12-28 16:56:15
description: decode field by opcode
*/

// `include "D:/GitHub/openx86/w80386dx/rtl/definition.h"
interface decode_interface (
    logic        opcode_MOV_reg_to_reg_mem,
    logic        opcode_MOV_reg_mem_to_reg,
    logic        opcode_MOV_imm_to_reg_mem,
    logic        opcode_MOV_imm_to_reg_short,
    logic        opcode_MOV_mem_to_acc,
    logic        opcode_MOV_acc_to_mem,
    logic        opcode_MOV_reg_mem_to_sreg,
    logic        opcode_MOV_sreg_to_reg_mem,
    logic        opcode_MOVSX,
    logic        opcode_MOVZX,
    logic        opcode_PUSH_reg_mem,
    logic        opcode_PUSH_reg_short,
    logic        opcode_PUSH_sreg_2,
    logic        opcode_PUSH_sreg_3,
    logic        opcode_PUSH_imm,
    logic        opcode_PUSH_all,
    logic        opcode_POP_reg_mem,
    logic        opcode_POP_reg_short,
    logic        opcode_POP_sreg_2,
    logic        opcode_POP_sreg_3,
    logic        opcode_POP_all,
    logic        opcode_XCHG_reg_mem_with_reg,
    logic        opcode_XCHG_reg_with_acc_short,
    logic        opcode_IN_port_fixed,
    logic        opcode_IN_port_variable,
    logic        opcode_OUT_port_fixed,
    logic        opcode_OUT_port_variable,
    logic        opcode_LEA_load_ea_to_reg,
    logic        opcode_LDS_load_ptr_to_DS,
    logic        opcode_LES_load_ptr_to_ES,
    logic        opcode_LFS_load_ptr_to_FS,
    logic        opcode_LGS_load_ptr_to_GS,
    logic        opcode_LSS_load_ptr_to_SS,
    logic        opcode_CLC_clear_carry_flag,
    logic        opcode_CLD_clear_direction_flag,
    logic        opcode_CLI_clear_interrupt_enable_flag,
    logic        opcode_CLTS_clear_task_switched_flag,
    logic        opcode_CMC_complement_carry_flag,
    logic        opcode_LAHF_load_ah_into_flag,
    logic        opcode_POPF_pop_flags,
    logic        opcode_PUSHF_push_flags,
    logic        opcode_SAHF_store_ah_into_flag,
    logic        opcode_STC_set_carry_flag,
    logic        opcode_STD_set_direction_flag,
    logic        opcode_STI_set_interrupt_enable_flag,
    logic        opcode_ADD_reg_to_mem,
    logic        opcode_ADD_mem_to_reg,
    logic        opcode_ADD_imm_to_reg_mem,
    logic        opcode_ADD_imm_to_acc,
    logic        opcode_ADC_reg_to_mem,
    logic        opcode_ADC_mem_to_reg,
    logic        opcode_ADC_imm_to_reg_mem,
    logic        opcode_ADC_imm_to_acc,
    logic        opcode_INC_reg_mem,
    logic        opcode_INC_reg,
    logic        opcode_SUB_reg_to_mem,
    logic        opcode_SUB_mem_to_reg,
    logic        opcode_SUB_imm_to_reg_mem,
    logic        opcode_SUB_imm_to_acc,
    logic        opcode_SBB_reg_to_mem,
    logic        opcode_SBB_mem_to_reg,
    logic        opcode_SBB_imm_to_reg_mem,
    logic        opcode_SBB_imm_to_acc,
    logic        opcode_DEC_reg_mem,
    logic        opcode_DEC_reg,
    logic        opcode_CMP_mem_with_reg,
    logic        opcode_CMP_reg_with_mem,
    logic        opcode_CMP_imm_with_reg_mem,
    logic        opcode_CMP_imm_with_acc,
    logic        opcode_NEG_change_sign,
    logic        opcode_AAA,
    logic        opcode_AAS,
    logic        opcode_DAA,
    logic        opcode_DAS,
    logic        opcode_MUL_acc_with_reg_mem,
    logic        opcode_IMUL_acc_with_reg_mem,
    logic        opcode_IMUL_reg_with_reg_mem,
    logic        opcode_IMUL_reg_mem_with_imm_to_reg,
    logic        opcode_DIV_acc_by_reg_mem,
    logic        opcode_IDIV_acc_by_reg_mem,
    logic        opcode_AAD,
    logic        opcode_AAM,
    logic        opcode_CBW,
    logic        opcode_CWD,
    logic        opcode_ROL_reg_mem_by_1,
    logic        opcode_ROL_reg_mem_by_CL,
    logic        opcode_ROL_reg_mem_by_imm,
    logic        opcode_ROR_reg_mem_by_1,
    logic        opcode_ROR_reg_mem_by_CL,
    logic        opcode_ROR_reg_mem_by_imm,
    logic        opcode_SHL_reg_mem_by_1,
    logic        opcode_SHL_reg_mem_by_CL,
    logic        opcode_SHL_reg_mem_by_imm,
    logic        opcode_SAR_reg_mem_by_1,
    logic        opcode_SAR_reg_mem_by_CL,
    logic        opcode_SAR_reg_mem_by_imm,
    logic        opcode_SHR_reg_mem_by_1,
    logic        opcode_SHR_reg_mem_by_CL,
    logic        opcode_SHR_reg_mem_by_imm,
    logic        opcode_RCL_reg_mem_by_1,
    logic        opcode_RCL_reg_mem_by_CL,
    logic        opcode_RCL_reg_mem_by_imm,
    logic        opcode_RCR_reg_mem_by_1,
    logic        opcode_RCR_reg_mem_by_CL,
    logic        opcode_RCR_reg_mem_by_imm,
    logic        opcode_SHLD_reg_mem_by_imm,
    logic        opcode_SHLD_reg_mem_by_CL,
    logic        opcode_SHRD_reg_mem_by_imm,
    logic        opcode_SHRD_reg_mem_by_CL,
    logic        opcode_AND_reg_to_mem,
    logic        opcode_AND_mem_to_reg,
    logic        opcode_AND_imm_to_reg_mem,
    logic        opcode_AND_imm_to_acc,
    logic        opcode_TEST_reg_mem_and_reg,
    logic        opcode_TEST_imm_to_reg_mem,
    logic        opcode_TEST_imm_to_acc,
    logic        opcode_OR_reg_to_mem,
    logic        opcode_OR_mem_to_reg,
    logic        opcode_OR_imm_to_reg_mem,
    logic        opcode_OR_imm_to_acc,
    logic        opcode_XOR_reg_to_mem,
    logic        opcode_XOR_mem_to_reg,
    logic        opcode_XOR_imm_to_reg_mem,
    logic        opcode_XOR_imm_to_acc,
    logic        opcode_NOT,
    logic        opcode_CMPS,
    logic        opcode_INS,
    logic        opcode_LODS,
    logic        opcode_MOVS,
    logic        opcode_OUTS,
    logic        opcode_SCAS,
    logic        opcode_STOS,
    logic        opcode_XLAT,
    logic        opcode_REPE,
    logic        opcode_REPNE,
    logic        opcode_BSF,
    logic        opcode_BSR,
    logic        opcode_BT_reg_mem_with_imm,
    logic        opcode_BT_reg_mem_with_reg,
    logic        opcode_BTC_reg_mem_with_imm,
    logic        opcode_BTC_reg_mem_with_reg,
    logic        opcode_BTR_reg_mem_with_imm,
    logic        opcode_BTR_reg_mem_with_reg,
    logic        opcode_BTS_reg_mem_with_imm,
    logic        opcode_BTS_reg_mem_with_reg,
    logic        opcode_CALL_direct_within_segment,
    logic        opcode_CALL_indirect_within_segment,
    logic        opcode_CALL_direct_intersegment,
    logic        opcode_CALL_indirect_intersegment,
    logic        opcode_JMP_short,
    logic        opcode_JMP_direct_within_segment,
    logic        opcode_JMP_indirect_within_segment,
    logic        opcode_JMP_direct_intersegment,
    logic        opcode_JMP_indirect_intersegment,
    logic        opcode_RET_within_segment,
    logic        opcode_RET_within_segment_adding_imm_to_SP,
    logic        opcode_RET_intersegment,
    logic        opcode_RET_intersegment_adding_imm_to_SP,
    logic        opcode_JO_8bit_disp,
    logic        opcode_JO_full_disp,
    logic        opcode_JNO_8bit_disp,
    logic        opcode_JNO_full_disp,
    logic        opcode_JB_8bit_disp,
    logic        opcode_JB_full_disp,
    logic        opcode_JNB_8bit_disp,
    logic        opcode_JNB_full_disp,
    logic        opcode_JE_8bit_disp,
    logic        opcode_JE_full_disp,
    logic        opcode_JNE_8bit_disp,
    logic        opcode_JNE_full_disp,
    logic        opcode_JBE_8bit_disp,
    logic        opcode_JBE_full_disp,
    logic        opcode_JNBE_8bit_disp,
    logic        opcode_JNBE_full_disp,
    logic        opcode_JS_8bit_disp,
    logic        opcode_JS_full_disp,
    logic        opcode_JNS_8bit_disp,
    logic        opcode_JNS_full_disp,
    logic        opcode_JP_8bit_disp,
    logic        opcode_JP_full_disp,
    logic        opcode_JNP_8bit_disp,
    logic        opcode_JNP_full_disp,
    logic        opcode_JL_8bit_disp,
    logic        opcode_JL_full_disp,
    logic        opcode_JNL_8bit_disp,
    logic        opcode_JNL_full_disp,
    logic        opcode_JLE_8bit_disp,
    logic        opcode_JLE_full_disp,
    logic        opcode_JNLE_8bit_disp,
    logic        opcode_JNLE_full_disp,
    logic        opcode_JCXZ,
    logic        opcode_LOOP,
    logic        opcode_LOOPZ,
    logic        opcode_LOOPNZ,
    logic        opcode_SETO,
    logic        opcode_SETNO,
    logic        opcode_SETB,
    logic        opcode_SETNB,
    logic        opcode_SETE,
    logic        opcode_SETNE,
    logic        opcode_SETBE,
    logic        opcode_SETNBE,
    logic        opcode_SETS,
    logic        opcode_SETNS,
    logic        opcode_SETP,
    logic        opcode_SETNP,
    logic        opcode_SETL,
    logic        opcode_SETNL,
    logic        opcode_SETLE,
    logic        opcode_SETNLE,
    logic        opcode_ENTER,
    logic        opcode_LEAVE,
    logic        opcode_INT_type_3,
    logic        opcode_INT_type_specified,
    logic        opcode_INTO,
    logic        opcode_BOUND,
    logic        opcode_IRET,
    logic        opcode_HLT,
    logic        opcode_MOV_CR0_CR2_CR3_from_reg,
    logic        opcode_MOV_reg_from_CR0_3,
    logic        opcode_MOV_DR0_7_from_reg,
    logic        opcode_MOV_reg_from_DR0_7,
    logic        opcode_MOV_TR6_7_from_reg,
    logic        opcode_MOV_reg_from_TR6_7,
    logic        opcode_NOP,
    logic        opcode_WAIT,
    logic        opcode_processor_extension_escape,
    logic        opcode_prefix_address_size,
    logic        opcode_prefix_bus_lock,
    logic        opcode_prefix_operand_size,
    logic        opcode_prefix_segment_override_CS,
    logic        opcode_prefix_segment_override_DS,
    logic        opcode_prefix_segment_override_ES,
    logic        opcode_prefix_segment_override_FS,
    logic        opcode_prefix_segment_override_GS,
    logic        opcode_prefix_segment_override_SS,
    logic        opcode_ARPL,
    logic        opcode_LAR,
    logic        opcode_LGDT,
    logic        opcode_LIDT,
    logic        opcode_LLDT,
    logic        opcode_LMSW,
    logic        opcode_LSL,
    logic        opcode_LTR,
    logic        opcode_SGDT,
    logic        opcode_SIDT,
    logic        opcode_SLDT,
    logic        opcode_SMSW,
    logic        opcode_STR,
    logic        opcode_VERR,
    logic        opcode_VERW
);

modport opcode_input (
    input  logic        opcode_MOV_reg_to_reg_mem,
    input  logic        opcode_MOV_reg_mem_to_reg,
    input  logic        opcode_MOV_imm_to_reg_mem,
    input  logic        opcode_MOV_imm_to_reg_short,
    input  logic        opcode_MOV_mem_to_acc,
    input  logic        opcode_MOV_acc_to_mem,
    input  logic        opcode_MOV_reg_mem_to_sreg,
    input  logic        opcode_MOV_sreg_to_reg_mem,
    input  logic        opcode_MOVSX,
    input  logic        opcode_MOVZX,
    input  logic        opcode_PUSH_reg_mem,
    input  logic        opcode_PUSH_reg_short,
    input  logic        opcode_PUSH_sreg_2,
    input  logic        opcode_PUSH_sreg_3,
    input  logic        opcode_PUSH_imm,
    input  logic        opcode_PUSH_all,
    input  logic        opcode_POP_reg_mem,
    input  logic        opcode_POP_reg_short,
    input  logic        opcode_POP_sreg_2,
    input  logic        opcode_POP_sreg_3,
    input  logic        opcode_POP_all,
    input  logic        opcode_XCHG_reg_mem_with_reg,
    input  logic        opcode_XCHG_reg_with_acc_short,
    input  logic        opcode_IN_port_fixed,
    input  logic        opcode_IN_port_variable,
    input  logic        opcode_OUT_port_fixed,
    input  logic        opcode_OUT_port_variable,
    input  logic        opcode_LEA_load_ea_to_reg,
    input  logic        opcode_LDS_load_ptr_to_DS,
    input  logic        opcode_LES_load_ptr_to_ES,
    input  logic        opcode_LFS_load_ptr_to_FS,
    input  logic        opcode_LGS_load_ptr_to_GS,
    input  logic        opcode_LSS_load_ptr_to_SS,
    input  logic        opcode_CLC_clear_carry_flag,
    input  logic        opcode_CLD_clear_direction_flag,
    input  logic        opcode_CLI_clear_interrupt_enable_flag,
    input  logic        opcode_CLTS_clear_task_switched_flag,
    input  logic        opcode_CMC_complement_carry_flag,
    input  logic        opcode_LAHF_load_ah_into_flag,
    input  logic        opcode_POPF_pop_flags,
    input  logic        opcode_PUSHF_push_flags,
    input  logic        opcode_SAHF_store_ah_into_flag,
    input  logic        opcode_STC_set_carry_flag,
    input  logic        opcode_STD_set_direction_flag,
    input  logic        opcode_STI_set_interrupt_enable_flag,
    input  logic        opcode_ADD_reg_to_mem,
    input  logic        opcode_ADD_mem_to_reg,
    input  logic        opcode_ADD_imm_to_reg_mem,
    input  logic        opcode_ADD_imm_to_acc,
    input  logic        opcode_ADC_reg_to_mem,
    input  logic        opcode_ADC_mem_to_reg,
    input  logic        opcode_ADC_imm_to_reg_mem,
    input  logic        opcode_ADC_imm_to_acc,
    input  logic        opcode_INC_reg_mem,
    input  logic        opcode_INC_reg,
    input  logic        opcode_SUB_reg_to_mem,
    input  logic        opcode_SUB_mem_to_reg,
    input  logic        opcode_SUB_imm_to_reg_mem,
    input  logic        opcode_SUB_imm_to_acc,
    input  logic        opcode_SBB_reg_to_mem,
    input  logic        opcode_SBB_mem_to_reg,
    input  logic        opcode_SBB_imm_to_reg_mem,
    input  logic        opcode_SBB_imm_to_acc,
    input  logic        opcode_DEC_reg_mem,
    input  logic        opcode_DEC_reg,
    input  logic        opcode_CMP_mem_with_reg,
    input  logic        opcode_CMP_reg_with_mem,
    input  logic        opcode_CMP_imm_with_reg_mem,
    input  logic        opcode_CMP_imm_with_acc,
    input  logic        opcode_NEG_change_sign,
    input  logic        opcode_AAA,
    input  logic        opcode_AAS,
    input  logic        opcode_DAA,
    input  logic        opcode_DAS,
    input  logic        opcode_MUL_acc_with_reg_mem,
    input  logic        opcode_IMUL_acc_with_reg_mem,
    input  logic        opcode_IMUL_reg_with_reg_mem,
    input  logic        opcode_IMUL_reg_mem_with_imm_to_reg,
    input  logic        opcode_DIV_acc_by_reg_mem,
    input  logic        opcode_IDIV_acc_by_reg_mem,
    input  logic        opcode_AAD,
    input  logic        opcode_AAM,
    input  logic        opcode_CBW,
    input  logic        opcode_CWD,
    input  logic        opcode_ROL_reg_mem_by_1,
    input  logic        opcode_ROL_reg_mem_by_CL,
    input  logic        opcode_ROL_reg_mem_by_imm,
    input  logic        opcode_ROR_reg_mem_by_1,
    input  logic        opcode_ROR_reg_mem_by_CL,
    input  logic        opcode_ROR_reg_mem_by_imm,
    input  logic        opcode_SHL_reg_mem_by_1,
    input  logic        opcode_SHL_reg_mem_by_CL,
    input  logic        opcode_SHL_reg_mem_by_imm,
    input  logic        opcode_SAR_reg_mem_by_1,
    input  logic        opcode_SAR_reg_mem_by_CL,
    input  logic        opcode_SAR_reg_mem_by_imm,
    input  logic        opcode_SHR_reg_mem_by_1,
    input  logic        opcode_SHR_reg_mem_by_CL,
    input  logic        opcode_SHR_reg_mem_by_imm,
    input  logic        opcode_RCL_reg_mem_by_1,
    input  logic        opcode_RCL_reg_mem_by_CL,
    input  logic        opcode_RCL_reg_mem_by_imm,
    input  logic        opcode_RCR_reg_mem_by_1,
    input  logic        opcode_RCR_reg_mem_by_CL,
    input  logic        opcode_RCR_reg_mem_by_imm,
    input  logic        opcode_SHLD_reg_mem_by_imm,
    input  logic        opcode_SHLD_reg_mem_by_CL,
    input  logic        opcode_SHRD_reg_mem_by_imm,
    input  logic        opcode_SHRD_reg_mem_by_CL,
    input  logic        opcode_AND_reg_to_mem,
    input  logic        opcode_AND_mem_to_reg,
    input  logic        opcode_AND_imm_to_reg_mem,
    input  logic        opcode_AND_imm_to_acc,
    input  logic        opcode_TEST_reg_mem_and_reg,
    input  logic        opcode_TEST_imm_to_reg_mem,
    input  logic        opcode_TEST_imm_to_acc,
    input  logic        opcode_OR_reg_to_mem,
    input  logic        opcode_OR_mem_to_reg,
    input  logic        opcode_OR_imm_to_reg_mem,
    input  logic        opcode_OR_imm_to_acc,
    input  logic        opcode_XOR_reg_to_mem,
    input  logic        opcode_XOR_mem_to_reg,
    input  logic        opcode_XOR_imm_to_reg_mem,
    input  logic        opcode_XOR_imm_to_acc,
    input  logic        opcode_NOT,
    input  logic        opcode_CMPS,
    input  logic        opcode_INS,
    input  logic        opcode_LODS,
    input  logic        opcode_MOVS,
    input  logic        opcode_OUTS,
    input  logic        opcode_SCAS,
    input  logic        opcode_STOS,
    input  logic        opcode_XLAT,
    input  logic        opcode_REPE,
    input  logic        opcode_REPNE,
    input  logic        opcode_BSF,
    input  logic        opcode_BSR,
    input  logic        opcode_BT_reg_mem_with_imm,
    input  logic        opcode_BT_reg_mem_with_reg,
    input  logic        opcode_BTC_reg_mem_with_imm,
    input  logic        opcode_BTC_reg_mem_with_reg,
    input  logic        opcode_BTR_reg_mem_with_imm,
    input  logic        opcode_BTR_reg_mem_with_reg,
    input  logic        opcode_BTS_reg_mem_with_imm,
    input  logic        opcode_BTS_reg_mem_with_reg,
    input  logic        opcode_CALL_direct_within_segment,
    input  logic        opcode_CALL_indirect_within_segment,
    input  logic        opcode_CALL_direct_intersegment,
    input  logic        opcode_CALL_indirect_intersegment,
    input  logic        opcode_JMP_short,
    input  logic        opcode_JMP_direct_within_segment,
    input  logic        opcode_JMP_indirect_within_segment,
    input  logic        opcode_JMP_direct_intersegment,
    input  logic        opcode_JMP_indirect_intersegment,
    input  logic        opcode_RET_within_segment,
    input  logic        opcode_RET_within_segment_adding_imm_to_SP,
    input  logic        opcode_RET_intersegment,
    input  logic        opcode_RET_intersegment_adding_imm_to_SP,
    input  logic        opcode_JO_8bit_disp,
    input  logic        opcode_JO_full_disp,
    input  logic        opcode_JNO_8bit_disp,
    input  logic        opcode_JNO_full_disp,
    input  logic        opcode_JB_8bit_disp,
    input  logic        opcode_JB_full_disp,
    input  logic        opcode_JNB_8bit_disp,
    input  logic        opcode_JNB_full_disp,
    input  logic        opcode_JE_8bit_disp,
    input  logic        opcode_JE_full_disp,
    input  logic        opcode_JNE_8bit_disp,
    input  logic        opcode_JNE_full_disp,
    input  logic        opcode_JBE_8bit_disp,
    input  logic        opcode_JBE_full_disp,
    input  logic        opcode_JNBE_8bit_disp,
    input  logic        opcode_JNBE_full_disp,
    input  logic        opcode_JS_8bit_disp,
    input  logic        opcode_JS_full_disp,
    input  logic        opcode_JNS_8bit_disp,
    input  logic        opcode_JNS_full_disp,
    input  logic        opcode_JP_8bit_disp,
    input  logic        opcode_JP_full_disp,
    input  logic        opcode_JNP_8bit_disp,
    input  logic        opcode_JNP_full_disp,
    input  logic        opcode_JL_8bit_disp,
    input  logic        opcode_JL_full_disp,
    input  logic        opcode_JNL_8bit_disp,
    input  logic        opcode_JNL_full_disp,
    input  logic        opcode_JLE_8bit_disp,
    input  logic        opcode_JLE_full_disp,
    input  logic        opcode_JNLE_8bit_disp,
    input  logic        opcode_JNLE_full_disp,
    input  logic        opcode_JCXZ,
    input  logic        opcode_LOOP,
    input  logic        opcode_LOOPZ,
    input  logic        opcode_LOOPNZ,
    input  logic        opcode_SETO,
    input  logic        opcode_SETNO,
    input  logic        opcode_SETB,
    input  logic        opcode_SETNB,
    input  logic        opcode_SETE,
    input  logic        opcode_SETNE,
    input  logic        opcode_SETBE,
    input  logic        opcode_SETNBE,
    input  logic        opcode_SETS,
    input  logic        opcode_SETNS,
    input  logic        opcode_SETP,
    input  logic        opcode_SETNP,
    input  logic        opcode_SETL,
    input  logic        opcode_SETNL,
    input  logic        opcode_SETLE,
    input  logic        opcode_SETNLE,
    input  logic        opcode_ENTER,
    input  logic        opcode_LEAVE,
    input  logic        opcode_INT_type_3,
    input  logic        opcode_INT_type_specified,
    input  logic        opcode_INTO,
    input  logic        opcode_BOUND,
    input  logic        opcode_IRET,
    input  logic        opcode_HLT,
    input  logic        opcode_MOV_CR0_CR2_CR3_from_reg,
    input  logic        opcode_MOV_reg_from_CR0_3,
    input  logic        opcode_MOV_DR0_7_from_reg,
    input  logic        opcode_MOV_reg_from_DR0_7,
    input  logic        opcode_MOV_TR6_7_from_reg,
    input  logic        opcode_MOV_reg_from_TR6_7,
    input  logic        opcode_NOP,
    input  logic        opcode_WAIT,
    input  logic        opcode_processor_extension_escape,
    input  logic        opcode_prefix_address_size,
    input  logic        opcode_prefix_bus_lock,
    input  logic        opcode_prefix_operand_size,
    input  logic        opcode_prefix_segment_override_CS,
    input  logic        opcode_prefix_segment_override_DS,
    input  logic        opcode_prefix_segment_override_ES,
    input  logic        opcode_prefix_segment_override_FS,
    input  logic        opcode_prefix_segment_override_GS,
    input  logic        opcode_prefix_segment_override_SS,
    input  logic        opcode_ARPL,
    input  logic        opcode_LAR,
    input  logic        opcode_LGDT,
    input  logic        opcode_LIDT,
    input  logic        opcode_LLDT,
    input  logic        opcode_LMSW,
    input  logic        opcode_LSL,
    input  logic        opcode_LTR,
    input  logic        opcode_SGDT,
    input  logic        opcode_SIDT,
    input  logic        opcode_SLDT,
    input  logic        opcode_SMSW,
    input  logic        opcode_STR,
    input  logic        opcode_VERR,
    input  logic        opcode_VERW
);

modport opcode_output (
    output logic        opcode_MOV_reg_to_reg_mem,
    output logic        opcode_MOV_reg_mem_to_reg,
    output logic        opcode_MOV_imm_to_reg_mem,
    output logic        opcode_MOV_imm_to_reg_short,
    output logic        opcode_MOV_mem_to_acc,
    output logic        opcode_MOV_acc_to_mem,
    output logic        opcode_MOV_reg_mem_to_sreg,
    output logic        opcode_MOV_sreg_to_reg_mem,
    output logic        opcode_MOVSX,
    output logic        opcode_MOVZX,
    output logic        opcode_PUSH_reg_mem,
    output logic        opcode_PUSH_reg_short,
    output logic        opcode_PUSH_sreg_2,
    output logic        opcode_PUSH_sreg_3,
    output logic        opcode_PUSH_imm,
    output logic        opcode_PUSH_all,
    output logic        opcode_POP_reg_mem,
    output logic        opcode_POP_reg_short,
    output logic        opcode_POP_sreg_2,
    output logic        opcode_POP_sreg_3,
    output logic        opcode_POP_all,
    output logic        opcode_XCHG_reg_mem_with_reg,
    output logic        opcode_XCHG_reg_with_acc_short,
    output logic        opcode_IN_port_fixed,
    output logic        opcode_IN_port_variable,
    output logic        opcode_OUT_port_fixed,
    output logic        opcode_OUT_port_variable,
    output logic        opcode_LEA_load_ea_to_reg,
    output logic        opcode_LDS_load_ptr_to_DS,
    output logic        opcode_LES_load_ptr_to_ES,
    output logic        opcode_LFS_load_ptr_to_FS,
    output logic        opcode_LGS_load_ptr_to_GS,
    output logic        opcode_LSS_load_ptr_to_SS,
    output logic        opcode_CLC_clear_carry_flag,
    output logic        opcode_CLD_clear_direction_flag,
    output logic        opcode_CLI_clear_interrupt_enable_flag,
    output logic        opcode_CLTS_clear_task_switched_flag,
    output logic        opcode_CMC_complement_carry_flag,
    output logic        opcode_LAHF_load_ah_into_flag,
    output logic        opcode_POPF_pop_flags,
    output logic        opcode_PUSHF_push_flags,
    output logic        opcode_SAHF_store_ah_into_flag,
    output logic        opcode_STC_set_carry_flag,
    output logic        opcode_STD_set_direction_flag,
    output logic        opcode_STI_set_interrupt_enable_flag,
    output logic        opcode_ADD_reg_to_mem,
    output logic        opcode_ADD_mem_to_reg,
    output logic        opcode_ADD_imm_to_reg_mem,
    output logic        opcode_ADD_imm_to_acc,
    output logic        opcode_ADC_reg_to_mem,
    output logic        opcode_ADC_mem_to_reg,
    output logic        opcode_ADC_imm_to_reg_mem,
    output logic        opcode_ADC_imm_to_acc,
    output logic        opcode_INC_reg_mem,
    output logic        opcode_INC_reg,
    output logic        opcode_SUB_reg_to_mem,
    output logic        opcode_SUB_mem_to_reg,
    output logic        opcode_SUB_imm_to_reg_mem,
    output logic        opcode_SUB_imm_to_acc,
    output logic        opcode_SBB_reg_to_mem,
    output logic        opcode_SBB_mem_to_reg,
    output logic        opcode_SBB_imm_to_reg_mem,
    output logic        opcode_SBB_imm_to_acc,
    output logic        opcode_DEC_reg_mem,
    output logic        opcode_DEC_reg,
    output logic        opcode_CMP_mem_with_reg,
    output logic        opcode_CMP_reg_with_mem,
    output logic        opcode_CMP_imm_with_reg_mem,
    output logic        opcode_CMP_imm_with_acc,
    output logic        opcode_NEG_change_sign,
    output logic        opcode_AAA,
    output logic        opcode_AAS,
    output logic        opcode_DAA,
    output logic        opcode_DAS,
    output logic        opcode_MUL_acc_with_reg_mem,
    output logic        opcode_IMUL_acc_with_reg_mem,
    output logic        opcode_IMUL_reg_with_reg_mem,
    output logic        opcode_IMUL_reg_mem_with_imm_to_reg,
    output logic        opcode_DIV_acc_by_reg_mem,
    output logic        opcode_IDIV_acc_by_reg_mem,
    output logic        opcode_AAD,
    output logic        opcode_AAM,
    output logic        opcode_CBW,
    output logic        opcode_CWD,
    output logic        opcode_ROL_reg_mem_by_1,
    output logic        opcode_ROL_reg_mem_by_CL,
    output logic        opcode_ROL_reg_mem_by_imm,
    output logic        opcode_ROR_reg_mem_by_1,
    output logic        opcode_ROR_reg_mem_by_CL,
    output logic        opcode_ROR_reg_mem_by_imm,
    output logic        opcode_SHL_reg_mem_by_1,
    output logic        opcode_SHL_reg_mem_by_CL,
    output logic        opcode_SHL_reg_mem_by_imm,
    output logic        opcode_SAR_reg_mem_by_1,
    output logic        opcode_SAR_reg_mem_by_CL,
    output logic        opcode_SAR_reg_mem_by_imm,
    output logic        opcode_SHR_reg_mem_by_1,
    output logic        opcode_SHR_reg_mem_by_CL,
    output logic        opcode_SHR_reg_mem_by_imm,
    output logic        opcode_RCL_reg_mem_by_1,
    output logic        opcode_RCL_reg_mem_by_CL,
    output logic        opcode_RCL_reg_mem_by_imm,
    output logic        opcode_RCR_reg_mem_by_1,
    output logic        opcode_RCR_reg_mem_by_CL,
    output logic        opcode_RCR_reg_mem_by_imm,
    output logic        opcode_SHLD_reg_mem_by_imm,
    output logic        opcode_SHLD_reg_mem_by_CL,
    output logic        opcode_SHRD_reg_mem_by_imm,
    output logic        opcode_SHRD_reg_mem_by_CL,
    output logic        opcode_AND_reg_to_mem,
    output logic        opcode_AND_mem_to_reg,
    output logic        opcode_AND_imm_to_reg_mem,
    output logic        opcode_AND_imm_to_acc,
    output logic        opcode_TEST_reg_mem_and_reg,
    output logic        opcode_TEST_imm_to_reg_mem,
    output logic        opcode_TEST_imm_to_acc,
    output logic        opcode_OR_reg_to_mem,
    output logic        opcode_OR_mem_to_reg,
    output logic        opcode_OR_imm_to_reg_mem,
    output logic        opcode_OR_imm_to_acc,
    output logic        opcode_XOR_reg_to_mem,
    output logic        opcode_XOR_mem_to_reg,
    output logic        opcode_XOR_imm_to_reg_mem,
    output logic        opcode_XOR_imm_to_acc,
    output logic        opcode_NOT,
    output logic        opcode_CMPS,
    output logic        opcode_INS,
    output logic        opcode_LODS,
    output logic        opcode_MOVS,
    output logic        opcode_OUTS,
    output logic        opcode_SCAS,
    output logic        opcode_STOS,
    output logic        opcode_XLAT,
    output logic        opcode_REPE,
    output logic        opcode_REPNE,
    output logic        opcode_BSF,
    output logic        opcode_BSR,
    output logic        opcode_BT_reg_mem_with_imm,
    output logic        opcode_BT_reg_mem_with_reg,
    output logic        opcode_BTC_reg_mem_with_imm,
    output logic        opcode_BTC_reg_mem_with_reg,
    output logic        opcode_BTR_reg_mem_with_imm,
    output logic        opcode_BTR_reg_mem_with_reg,
    output logic        opcode_BTS_reg_mem_with_imm,
    output logic        opcode_BTS_reg_mem_with_reg,
    output logic        opcode_CALL_direct_within_segment,
    output logic        opcode_CALL_indirect_within_segment,
    output logic        opcode_CALL_direct_intersegment,
    output logic        opcode_CALL_indirect_intersegment,
    output logic        opcode_JMP_short,
    output logic        opcode_JMP_direct_within_segment,
    output logic        opcode_JMP_indirect_within_segment,
    output logic        opcode_JMP_direct_intersegment,
    output logic        opcode_JMP_indirect_intersegment,
    output logic        opcode_RET_within_segment,
    output logic        opcode_RET_within_segment_adding_imm_to_SP,
    output logic        opcode_RET_intersegment,
    output logic        opcode_RET_intersegment_adding_imm_to_SP,
    output logic        opcode_JO_8bit_disp,
    output logic        opcode_JO_full_disp,
    output logic        opcode_JNO_8bit_disp,
    output logic        opcode_JNO_full_disp,
    output logic        opcode_JB_8bit_disp,
    output logic        opcode_JB_full_disp,
    output logic        opcode_JNB_8bit_disp,
    output logic        opcode_JNB_full_disp,
    output logic        opcode_JE_8bit_disp,
    output logic        opcode_JE_full_disp,
    output logic        opcode_JNE_8bit_disp,
    output logic        opcode_JNE_full_disp,
    output logic        opcode_JBE_8bit_disp,
    output logic        opcode_JBE_full_disp,
    output logic        opcode_JNBE_8bit_disp,
    output logic        opcode_JNBE_full_disp,
    output logic        opcode_JS_8bit_disp,
    output logic        opcode_JS_full_disp,
    output logic        opcode_JNS_8bit_disp,
    output logic        opcode_JNS_full_disp,
    output logic        opcode_JP_8bit_disp,
    output logic        opcode_JP_full_disp,
    output logic        opcode_JNP_8bit_disp,
    output logic        opcode_JNP_full_disp,
    output logic        opcode_JL_8bit_disp,
    output logic        opcode_JL_full_disp,
    output logic        opcode_JNL_8bit_disp,
    output logic        opcode_JNL_full_disp,
    output logic        opcode_JLE_8bit_disp,
    output logic        opcode_JLE_full_disp,
    output logic        opcode_JNLE_8bit_disp,
    output logic        opcode_JNLE_full_disp,
    output logic        opcode_JCXZ,
    output logic        opcode_LOOP,
    output logic        opcode_LOOPZ,
    output logic        opcode_LOOPNZ,
    output logic        opcode_SETO,
    output logic        opcode_SETNO,
    output logic        opcode_SETB,
    output logic        opcode_SETNB,
    output logic        opcode_SETE,
    output logic        opcode_SETNE,
    output logic        opcode_SETBE,
    output logic        opcode_SETNBE,
    output logic        opcode_SETS,
    output logic        opcode_SETNS,
    output logic        opcode_SETP,
    output logic        opcode_SETNP,
    output logic        opcode_SETL,
    output logic        opcode_SETNL,
    output logic        opcode_SETLE,
    output logic        opcode_SETNLE,
    output logic        opcode_ENTER,
    output logic        opcode_LEAVE,
    output logic        opcode_INT_type_3,
    output logic        opcode_INT_type_specified,
    output logic        opcode_INTO,
    output logic        opcode_BOUND,
    output logic        opcode_IRET,
    output logic        opcode_HLT,
    output logic        opcode_MOV_CR0_CR2_CR3_from_reg,
    output logic        opcode_MOV_reg_from_CR0_3,
    output logic        opcode_MOV_DR0_7_from_reg,
    output logic        opcode_MOV_reg_from_DR0_7,
    output logic        opcode_MOV_TR6_7_from_reg,
    output logic        opcode_MOV_reg_from_TR6_7,
    output logic        opcode_NOP,
    output logic        opcode_WAIT,
    output logic        opcode_processor_extension_escape,
    output logic        opcode_prefix_address_size,
    output logic        opcode_prefix_bus_lock,
    output logic        opcode_prefix_operand_size,
    output logic        opcode_prefix_segment_override_CS,
    output logic        opcode_prefix_segment_override_DS,
    output logic        opcode_prefix_segment_override_ES,
    output logic        opcode_prefix_segment_override_FS,
    output logic        opcode_prefix_segment_override_GS,
    output logic        opcode_prefix_segment_override_SS,
    output logic        opcode_ARPL,
    output logic        opcode_LAR,
    output logic        opcode_LGDT,
    output logic        opcode_LIDT,
    output logic        opcode_LLDT,
    output logic        opcode_LMSW,
    output logic        opcode_LSL,
    output logic        opcode_LTR,
    output logic        opcode_SGDT,
    output logic        opcode_SIDT,
    output logic        opcode_SLDT,
    output logic        opcode_SMSW,
    output logic        opcode_STR,
    output logic        opcode_VERR,
    output logic        opcode_VERW
);

endinterface
